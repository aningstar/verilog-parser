module abc (id3, id4);

    input id3;
    output id4;

    reg signed a,b,c;
    reg a,b,c;
    reg scalared a,b,c;
    reg vectored a,b,c;
    reg [7:0] Q [0:3][0:15];
    reg signed [7:0] d1, d2;
    integer i, j;
    real r1, r2;
    real r1, r2;
    reg signed clock = 0, reset = 1;

endmodule
