module abc (id3, id4);
input signed [2:WORD] id3;
output  signed id4;

endmodule
