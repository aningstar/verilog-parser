module abc (id3, id4);

a = array1[1][2];

endmodule
