module abc (id3, id4);
    function automatic [63:0] factorial (input reg [31:0] n,t,r);
    endfunction

    function real multiply;
        input a, b;
    endfunction

    function Parity_Calc_Func;
         input [31:0] addr;
    endfunction

endmodule
