module abc (id3, id4);

endmodule