module abc (id3, id4);
out = 32'b11;
out = 32'o11;
out = 32'd11;
out = 32'h11;
endmodule