module abc (id3, id4);
input [5:0] id3;
output [6:8] id4;
reg e, k, l;

endmodule