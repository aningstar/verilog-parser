module abc (id3, id4);

    input id3;
    output id4;

    a = array1[1][2];

endmodule
