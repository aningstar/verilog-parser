module abc (id3, id4);
input signed [5:0] id3;
output  signed id4;

endmodule
