//`timescale 1ns/10ps

module pulse_delay (in, out);

input in;
output out;

wire n1, n2, n3, n4, n5, n6, n7, n8, n9, n10;

   inv_1 invi1 ( .x(n1), .a(in) );
   inv_1 invi2 ( .x(n2), .a(n1) );
   inv_1 invi3 ( .x(n3), .a(n2) );
   inv_1 invi4 ( .x(n4), .a(n3) );
   inv_1 invi5 ( .x(n5), .a(n4) );
   inv_1 invi6 ( .x(n6), .a(n5) );
   inv_1 invi7 ( .x(n7), .a(n6) );
   inv_1 invi8 ( .x(n8), .a(n7) );
   inv_1 invi9 ( .x(n9), .a(n8) );
   inv_1 invi10 ( .x(n10), .a(n9) );
   inv_1 invi11 ( .x(out), .a(n10) );

endmodule

module C_gate2 (  in1, in2, out );

input  in1, in2;
output  out;


	adfull_1 U3 ( .s(), .co(out), .a(in1), .b(in2), .ci(out) );

endmodule


module mymux4 (  mux_sel, out, in );

input [0:3] in;
input [1:0] mux_sel;
output  out;

	mux4_1 U4 ( .x(out), .d0(in[0]), .d1(in[1]), .d2(in[2]), .d3(in[3]), .sl0(mux_sel[0]), .sl1(mux_sel[1]) );

// mux4_1 U4 ( .x(out), .d0(in[0]), .d1(in[2]), .d2(in[1]), .d3(in[3]), .sl0(mux_sel[0]), .sl1(mux_sel[1]) ); //

endmodule


module matched_delay32__0_85__1__1_38__1_77 (  in, out, mux_sel );

input  in;
input [1:0] mux_sel;
output  out;

wire n1, n2, n3, net1, net10, net11, net12, net13, net14, net15, net16,
	net17, net18, net19, net2, net20, net21, net22, net23, net24, net25, net26,
	net27, net28, net29, net3, net30, net31, net32, net4, net5, net6, net7,
	net8, net9;

/*
pavlos 14 - 7
to n3 na odhghsei ola ta shmata
oi kathisterhseis na eine logarithmikis klimakas
*/
	buf_1 U1 ( .x(n1), .a(in) );
	buf_4 U2 ( .x(n2), .a(n1) );
	buf_16 U3 ( .x(n3), .a(n2) );
	and2_1 and1 ( .x(net1), .a(n3), .b(n3) );
        and2_1 and2 ( .x(net2), .a(n3), .b(net1) );
        and2_1 and3 ( .x(net3), .a(n3), .b(net2) );
        and2_1 and4 ( .x(net4), .a(n3), .b(net3) );
	and2_1 and5 ( .x(net5), .a(n3), .b(net4) );
	and2_1 and6 ( .x(net6), .a(n3), .b(net5) );
	and2_1 and7 ( .x(net7), .a(n3), .b(net6) );
	and2_1 and8 ( .x(net8), .a(n3), .b(net7) );
	and2_1 and9 ( .x(net9), .a(n3), .b(net8) );
	and2_1 and10 ( .x(net10), .a(n3), .b(net9) );
	and2_1 and11 ( .x(net11), .a(n3), .b(net10) );
	and2_1 and12 ( .x(net12), .a(n3), .b(net11) );
	and2_1 and13 ( .x(net13), .a(n3), .b(net12) );
	and2_1 and14 ( .x(net14), .a(n3), .b(net13) );
	and2_1 and15 ( .x(net15), .a(n3), .b(net14) );
	and2_1 and16 ( .x(net16), .a(n3), .b(net15) );
	and2_1 and17 ( .x(net17), .a(n3), .b(net16) );
	and2_1 and18 ( .x(net18), .a(n3), .b(net17) );
	and2_1 and19 ( .x(net19), .a(n3), .b(net18) );
	and2_1 and20 ( .x(net20), .a(n3), .b(net19) );
	/*and2_1 and21 ( .x(net21), .a(n3), .b(net20) );
	and2_1 and22 ( .x(net22), .a(n3), .b(net21) );
	and2_1 and23 ( .x(net23), .a(n3), .b(net22) );
	and2_1 and24 ( .x(net24), .a(n3), .b(net23) );
	and2_1 and25 ( .x(net25), .a(n3), .b(net24) );
	and2_1 and26 ( .x(net26), .a(n3), .b(net25) );
	and2_1 and27 ( .x(net27), .a(n3), .b(net26) );
	and2_1 and28 ( .x(net28), .a(n3), .b(net27) );
	and2_1 and29 ( .x(net29), .a(n3), .b(net28) );
	and2_1 and30 ( .x(net30), .a(n3), .b(net29) );
	and2_1 and31 ( .x(net31), .a(n3), .b(net30) );
	and2_1 and32 ( .x(net32), .a(n3), .b(net31) );*/


// mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net4, net8, net16, net32}) );

//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net15, net18, net25, net32}) );

//mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net13, net16, net20, net25}) );//1,25 logarithmic

mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net3, net5, net10, net20}) );//2 logarithmic

endmodule


module lc_semi_dec_master (  rst, ri, ai, ro, ao, l );

input  rst, ri, ao;
output  ai, ro, l;

wire aoi1, lint, nl, nri, nro, nrst;

	assign ai = nl;

	inv_1 linvg ( .x(l), .a(nl) );
	inv_1 linvi ( .x(lint), .a(nl) );
	aoi23_1 maingate ( .x(nl), .a(aoi1), .b(nri), .c(nri), .d(ro), .e(ao) );
	inv_1 resetinv ( .x(nrst), .a(rst) );
	nand2_1 resetnand ( .x(aoi1), .a(nrst), .b(ai) );
	inv_1 riinv ( .x(nri), .a(ri) );
	aoi21_1 rogate ( .x(ro), .a(nro), .b(ao), .c(lint) );
	inv_1 roint ( .x(nro), .a(ro) );

endmodule


module lc_semi_dec_slave (  rst, ri, ai, ro, ao, l );

input  rst, ri, ao;
output  ai, ro, l;

wire aoi1, lint, nl, nri, nro;

wire nri_del, naoi1_del, aoi1_del;

//        pulse_delay pulsedel ( ri, nri_del );
//        inv_1 temp ( .x(ri_del), .a(nri_del) );
//        pulse_delay pulsedel2 ( ri_del, nri_del_del );

	assign ai = nl;

	// delay of feedback (left input) must match pulse delay (right input) of LHS AND //

	inv_1 linvg ( .x(l), .a(nl) );
	inv_1 linvi ( .x(lint), .a(nl) );

//	aoi23_1 maingate ( .x(nl), .a(aoi1), .b(nri_del), .c(nri_del_del), .d(ro), .e(ao) );
   	aoi23_1 maingate ( .x(nl), .a(aoi1), .b(nri), .c(nri), .d(ro), .e(ao) );

	nor2_1 resetnor ( .x(aoi1), .a(rst), .b(ai) );
	inv_1 riinv ( .x(nri), .a(ri) );
	aoi221_1 rogate ( .x(ro), .a(nro), .b(ao), .c(lint), .d(1'b1), .e(rst) );
	inv_1 roint ( .x(nro), .a(ro) );

endmodule


module controller_d32__0_85__1__1_38__1_77_r1_a2 (  reset, en1, en2, ri1,
	ai, ro, ao1, ao2, delay_mux_sel );

input  reset, ri1, ao1, ao2;
input [1:0] delay_mux_sel;
output  en1, en2, ai, ro;

wire ao_synchr, ax, ri_synchr, ri_synchr_delayed, rx;

	assign ri_synchr = ri1;

	C_gate2 cgate_ackouts ( .in1(ao1), .in2(ao2), .out(ao_synchr) );
	matched_delay32__0_85__1__1_38__1_77 delay ( .in(ri_synchr), .out(ri_synchr_delayed),
		.mux_sel(delay_mux_sel) );
	lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai),
		.ro(rx), .ao(ax), .l(en1) );
	lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(ao_synchr),
		.l(en2) );

endmodule


module matched_delay31__0_85__1__1_47__1_93 (  in, out, mux_sel );

input  in;
input [1:0] mux_sel;
output  out;

wire n1, n2, n3, net1, net10, net11, net12, net13, net14, net15, net16,
	net17, net18, net19, net2, net20, net21, net22, net23, net24, net25, net26,
	net27, net28, net29, net3, net30, net31, net4, net5, net6, net7, net8,
	net9;


	buf_1 U1 ( .x(n1), .a(in) );
	buf_4 U2 ( .x(n2), .a(n1) );
	buf_16 U3 ( .x(n3), .a(n2) );
	and2_1 and1 ( .x(net1), .a(n3), .b(n3) );
        and2_1 and2 ( .x(net2), .a(n3), .b(net1) );
        and2_1 and3 ( .x(net3), .a(n3), .b(net2) );
        and2_1 and4 ( .x(net4), .a(n3), .b(net3) );
	and2_1 and5 ( .x(net5), .a(n3), .b(net4) );
	and2_1 and6 ( .x(net6), .a(n3), .b(net5) );
	and2_1 and7 ( .x(net7), .a(n3), .b(net6) );
	and2_1 and8 ( .x(net8), .a(n3), .b(net7) );
	and2_1 and9 ( .x(net9), .a(n3), .b(net8) );
	and2_1 and10 ( .x(net10), .a(n3), .b(net9) );
	and2_1 and11 ( .x(net11), .a(n3), .b(net10) );
	and2_1 and12 ( .x(net12), .a(n3), .b(net11) );
	and2_1 and13 ( .x(net13), .a(n3), .b(net12) );
	and2_1 and14 ( .x(net14), .a(n3), .b(net13) );
	and2_1 and15 ( .x(net15), .a(n3), .b(net14) );
	and2_1 and16 ( .x(net16), .a(n3), .b(net15) );
	and2_1 and17 ( .x(net17), .a(n3), .b(net16) );
	and2_1 and18 ( .x(net18), .a(n3), .b(net17) );
	and2_1 and19 ( .x(net19), .a(n3), .b(net18) );
	and2_1 and20 ( .x(net20), .a(n3), .b(net19) );
	/*and2_1 and21 ( .x(net21), .a(n3), .b(net20) );
	and2_1 and22 ( .x(net22), .a(n3), .b(net21) );
	and2_1 and23 ( .x(net23), .a(n3), .b(net22) );
	and2_1 and24 ( .x(net24), .a(n3), .b(net23) );
	and2_1 and25 ( .x(net25), .a(n3), .b(net24) );
	and2_1 and26 ( .x(net26), .a(n3), .b(net25) );
	and2_1 and27 ( .x(net27), .a(n3), .b(net26) );
	and2_1 and28 ( .x(net28), .a(n3), .b(net27) );
	and2_1 and29 ( .x(net29), .a(n3), .b(net28) );
	and2_1 and30 ( .x(net30), .a(n3), .b(net29) );
	and2_1 and31 ( .x(net31), .a(n3), .b(net30) );*/


//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net4, net8, net16, net31}) );

//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net13, net15, net24, net31}) );

//      mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net13, net16, net20, net24}) );//1,25 logarithmic

mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net3, net5, net10, net20}) );//2 logarithmic

endmodule


module controller_d31__0_85__1__1_47__1_93_r2_a2 (  reset, en1, en2, ri1,
	ri2, ai, ro, ao1, ao2, delay_mux_sel );

input  reset, ri1, ri2, ao1, ao2;
input [1:0] delay_mux_sel;
output  en1, en2, ai, ro;

wire ao_synchr, ax, ri_synchr, ri_synchr_delayed, rx;


	C_gate2 cgate_ackouts ( .in1(ao1), .in2(ao2), .out(ao_synchr) );
	C_gate2 cgate_reqins ( .in1(ri1), .in2(ri2), .out(ri_synchr) );
	matched_delay31__0_85__1__1_47__1_93 delay ( .in(ri_synchr), .out(ri_synchr_delayed),
		.mux_sel(delay_mux_sel) );
	lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai),
		.ro(rx), .ao(ax), .l(en1) );
	lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(ao_synchr),
		.l(en2) );

endmodule


module matched_delay28__0_85__1__1_48__1_95 (  in, out, mux_sel );

input  in;
input [1:0] mux_sel;
output  out;

wire n1, n2, n3, net1, net10, net11, net12, net13, net14, net15, net16,
	net17, net18, net19, net2, net20, net21, net22, net23, net24, net25, net26,
	net27, net28, net3, net4, net5, net6, net7, net8, net9;


	buf_1 U1 ( .x(n1), .a(in) );
	buf_4 U2 ( .x(n2), .a(n1) );
	buf_16 U3 ( .x(n3), .a(n2) );
	and2_1 and1 ( .x(net1), .a(n3), .b(n3) );
        and2_1 and2 ( .x(net2), .a(n3), .b(net1) );
        and2_1 and3 ( .x(net3), .a(n3), .b(net2) );
	and2_1 and4 ( .x(net4), .a(n3), .b(net3) );
	and2_1 and5 ( .x(net5), .a(n3), .b(net4) );
	and2_1 and6 ( .x(net6), .a(n3), .b(net5) );
	and2_1 and7 ( .x(net7), .a(n3), .b(net6) );
	and2_1 and8 ( .x(net8), .a(n3), .b(net7) );
	and2_1 and9 ( .x(net9), .a(n3), .b(net8) );
	and2_1 and10 ( .x(net10), .a(n3), .b(net9) );
	and2_1 and11 ( .x(net11), .a(n3), .b(net10) );
	and2_1 and12 ( .x(net12), .a(n3), .b(net11) );
	and2_1 and13 ( .x(net13), .a(n3), .b(net12) );
	and2_1 and14 ( .x(net14), .a(n3), .b(net13) );
	and2_1 and15 ( .x(net15), .a(n3), .b(net14) );
	and2_1 and16 ( .x(net16), .a(n3), .b(net15) );
	and2_1 and17 ( .x(net17), .a(n3), .b(net16) );
	and2_1 and18 ( .x(net18), .a(n3), .b(net17) );
	and2_1 and19 ( .x(net19), .a(n3), .b(net18) );
	and2_1 and20 ( .x(net20), .a(n3), .b(net19) );
	/*and2_1 and21 ( .x(net21), .a(n3), .b(net20) );
	and2_1 and22 ( .x(net22), .a(n3), .b(net21) );
	and2_1 and23 ( .x(net23), .a(n3), .b(net22) );
	and2_1 and24 ( .x(net24), .a(n3), .b(net23) );
	and2_1 and25 ( .x(net25), .a(n3), .b(net24) );
	and2_1 and26 ( .x(net26), .a(n3), .b(net25) );
	and2_1 and27 ( .x(net27), .a(n3), .b(net26) );
	and2_1 and28 ( .x(net28), .a(n3), .b(net27) );*/


//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net3, net7, net14, net28}) );

//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net11, net14, net21, net28}) );

//mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net13, net16, net20, net25}) );//1,25 logarithmic

mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net3, net5, net10, net20}) );//2 logarithmic

endmodule


module controller_d28__0_85__1__1_48__1_95_r2_a2 (  reset, en1, en2, ri1,
	ri2, ai, ro, ao1, ao2, delay_mux_sel );

input  reset, ri1, ri2, ao1, ao2;
input [1:0] delay_mux_sel;
output  en1, en2, ai, ro;

wire ao_synchr, ax, ri_synchr, ri_synchr_delayed, rx;


	C_gate2 cgate_ackouts ( .in1(ao1), .in2(ao2), .out(ao_synchr) );
	C_gate2 cgate_reqins ( .in1(ri1), .in2(ri2), .out(ri_synchr) );
	matched_delay28__0_85__1__1_48__1_95 delay ( .in(ri_synchr), .out(ri_synchr_delayed),
		.mux_sel(delay_mux_sel) );
	lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai),
		.ro(rx), .ao(ax), .l(en1) );
	lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(ao_synchr),
		.l(en2) );

endmodule


module matched_delay6__0_85__1__1_18__1_36 (  in, out, mux_sel );

input  in;
input [1:0] mux_sel;
output  out;

wire n1, n2, net1, net2, net3, net4, net5, net6;


	buf_1 U1 ( .x(n1), .a(in) );
	buf_4 U2 ( .x(n2), .a(n1) );
	and2_1 and1 ( .x(net1), .a(n2), .b(n2) );
	and2_1 and2 ( .x(net2), .a(n2), .b(net1) );
	and2_1 and3 ( .x(net3), .a(n2), .b(net2) );
	and2_1 and4 ( .x(net4), .a(n2), .b(net3) );
	and2_1 and5 ( .x(net5), .a(n2), .b(net4) );
	and2_1 and6 ( .x(net6), .a(n2), .b(net5) );

//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net1, net2, net4, net6}) );

//	mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net4, net4, net5, net6}) );

//mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net3, net4, net5, net6}) );//1,25 logarithmic

mymux4 mux ( .mux_sel(mux_sel), .out(out), .in({ net1, net2, net4, net6}) );//2 logarithmic

endmodule


module controller_d6__0_85__1__1_18__1_36_r2_a1 (  reset, en1, en2, ri1,
	ri2, ai, ro, ao1, delay_mux_sel );

input  reset, ri1, ri2, ao1;
input [1:0] delay_mux_sel;
output  en1, en2, ai, ro;

wire ao_synchr, ax, ri_synchr, ri_synchr_delayed, rx;

	assign ao_synchr = ao1;

	C_gate2 cgate_reqins ( .in1(ri1), .in2(ri2), .out(ri_synchr) );
	matched_delay6__0_85__1__1_18__1_36 delay ( .in(ri_synchr), .out(ri_synchr_delayed),
		.mux_sel(delay_mux_sel) );
	lc_semi_dec_master master ( .rst(reset), .ri(ri_synchr_delayed), .ai(ai),
		.ro(rx), .ao(ax), .l(en1) );
	lc_semi_dec_slave slave ( .rst(reset), .ri(rx), .ai(ax), .ro(ro), .ao(ao_synchr),
		.l(en2) );

endmodule


module smlatnr_2 (  q, qb, d, sdi, se, g, rb, glob_g, sync_sel );

input  d, sdi, se, g, rb, glob_g, sync_sel;
output  q, qb;

wire data, enable;


	latnr_2 latch ( .q(q), .qb(qb), .rb(rb), .d(data), .g(enable) );
	mux2_1 mux_scan ( .x(data), .d0(d), .sl(se), .d1(sdi) );
	mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );

endmodule


module mlatnr_8 (  q, qb, d, g, rb, glob_g, sync_sel );

input  d, g, rb, glob_g, sync_sel;
output  q, qb;

wire enable;


	latnr_8 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
	mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );

endmodule


module smlatnr_1 (  q, qb, d, sdi, se, g, rb, glob_g, sync_sel );

input  d, sdi, se, g, rb, glob_g, sync_sel;
output  q, qb;

wire data, enable;


	latnr_1 latch ( .q(q), .qb(qb), .rb(rb), .d(data), .g(enable) );
	mux2_1 mux_scan ( .x(data), .d0(d), .sl(se), .d1(sdi) );
	mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );

endmodule


module mlatnr_4 (  q, qb, d, g, rb, glob_g, sync_sel );

input  d, g, rb, glob_g, sync_sel;
output  q, qb;

wire enable;


	latnr_4 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
	mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );

endmodule


module mlatnr_2 (  q, qb, d, g, rb, glob_g, sync_sel );

input  d, g, rb, glob_g, sync_sel;
output  q, qb;

wire enable;


	latnr_2 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
	mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );

endmodule


module mlatnr_1 (  q, qb, d, g, rb, glob_g, sync_sel );

input  d, g, rb, glob_g, sync_sel;
output  q, qb;

wire enable;


	latnr_1 latch ( .q(q), .qb(qb), .rb(rb), .d(d), .g(enable) );
	mux2_1 mux_sync ( .x(enable), .d0(glob_g), .sl(sync_sel), .d1(g) );

endmodule


module EX_DW01_add_32_5_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
	n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
	n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
	n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
	n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
	n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
	n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
	n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
	n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
	n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
	n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n49,
	n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
	n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
	n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
	n92, n93, n94, n95, n96, n97, n98, n99;


	exnor2_5 U10 ( .x(SUM[30]), .a(n167), .b(n181) );
	inv_2 U100 ( .x(n367), .a(n313) );
	nand2_0 U101 ( .x(n365), .a(A[0]), .b(B[0]) );
	oai22_1 U102 ( .x(n322), .a(n224), .b(n225), .c(n250), .d(n321) );
	inv_2 U103 ( .x(n250), .a(n311) );
	inv_2 U104 ( .x(n321), .a(n174) );
	inv_2 U107 ( .x(n173), .a(n322) );
	inv_2 U108 ( .x(n96), .a(n251) );
	nor2i_1 U109 ( .x(n94), .a(n95), .b(n96) );
	nor2_2 U11 ( .x(n111), .a(A[15]), .b(B[15]) );
	inv_2 U110 ( .x(n330), .a(n138) );
	nand2i_2 U111 ( .x(n202), .a(n330), .b(n331) );
	inv_2 U112 ( .x(n332), .a(n202) );
	inv_0 U113 ( .x(n136), .a(n243) );
	oai21_1 U114 ( .x(n200), .a(n136), .b(n332), .c(n135) );
	exnor2_1 U115 ( .x(SUM[16]), .a(n199), .b(n131) );
	inv_5 U116 ( .x(n199), .a(n129) );
	nor2i_0 U117 ( .x(n131), .a(n132), .b(n133) );
	exor2_1 U118 ( .x(SUM[17]), .a(n197), .b(n198) );
	nor2_0 U12 ( .x(n170), .a(A[4]), .b(B[4]) );
	nand2i_2 U120 ( .x(n193), .a(n341), .b(n109) );
	inv_2 U121 ( .x(n161), .a(n109) );
	nand2i_0 U122 ( .x(n347), .a(n121), .b(n161) );
	nand2_0 U123 ( .x(n348), .a(A[22]), .b(B[22]) );
	inv_2 U124 ( .x(n341), .a(n159) );
	inv_0 U125 ( .x(n233), .a(B[21]) );
	nand2i_2 U126 ( .x(n314), .a(A[22]), .b(n107) );
	nand2i_2 U127 ( .x(n300), .a(n121), .b(n159) );
	nand2i_2 U128 ( .x(n190), .a(n342), .b(n343) );
	inv_2 U129 ( .x(n355), .a(n266) );
	or3i_2 U130 ( .x(n266), .a(n159), .b(n234), .c(n121) );
	aoi21_1 U131 ( .x(n294), .a(n272), .b(n295), .c(n296) );
	oai31_1 U132 ( .x(n272), .a(n108), .b(n121), .c(n110), .d(n273) );
	nand2i_0 U133 ( .x(n295), .a(B[24]), .b(n232) );
	inv_2 U134 ( .x(n296), .a(n343) );
	inv_2 U135 ( .x(n353), .a(n272) );
	inv_2 U136 ( .x(n234), .a(B[23]) );
	nand2i_2 U137 ( .x(n360), .a(n342), .b(n354) );
	inv_2 U138 ( .x(n342), .a(n295) );
	inv_2 U139 ( .x(n232), .a(A[24]) );
	inv_1 U14 ( .x(n242), .a(n363) );
	inv_2 U140 ( .x(n354), .a(n267) );
	or3i_2 U141 ( .x(n267), .a(n159), .b(n235), .c(n121) );
	inv_2 U142 ( .x(n235), .a(A[23]) );
	inv_2 U143 ( .x(n93), .a(n83) );
	nand2_2 U144 ( .x(n116), .a(A[25]), .b(B[25]) );
	inv_2 U145 ( .x(n119), .a(n211) );
	nor2i_1 U146 ( .x(n117), .a(n118), .b(n119) );
	inv_2 U147 ( .x(n182), .a(n307) );
	exnor2_1 U148 ( .x(SUM[3]), .a(n182), .b(n117) );
	exor2_1 U149 ( .x(SUM[2]), .a(n122), .b(n124) );
	inv_0 U15 ( .x(n263), .a(B[15]) );
	exor2_1 U150 ( .x(SUM[6]), .a(n177), .b(n100) );
	oai21_1 U151 ( .x(n177), .a(n371), .b(n178), .c(n104) );
	nor2i_1 U152 ( .x(n100), .a(n101), .b(n102) );
	exor2_1 U153 ( .x(SUM[12]), .a(n204), .b(n140) );
	exor2_1 U154 ( .x(SUM[7]), .a(n176), .b(n97) );
	oai21_1 U155 ( .x(n176), .a(n102), .b(n325), .c(n101) );
	inv_0 U156 ( .x(n102), .a(n310) );
	inv_2 U157 ( .x(n325), .a(n177) );
	nor2i_1 U158 ( .x(n97), .a(n98), .b(n99) );
	inv_2 U159 ( .x(n99), .a(n287) );
	nand2i_2 U16 ( .x(n275), .a(n138), .b(n243) );
	exor2_1 U160 ( .x(n186), .a(B[27]), .b(A[27]) );
	exor2_1 U162 ( .x(n195), .a(A[20]), .b(B[20]) );
	exor2_1 U163 ( .x(SUM[14]), .a(n202), .b(n134) );
	exor2_1 U164 ( .x(SUM[10]), .a(n206), .b(n146) );
	nor2i_0 U165 ( .x(n103), .a(n104), .b(n371) );
	inv_2 U166 ( .x(n323), .a(n179) );
	aoai211_1 U167 ( .x(n324), .a(n217), .b(n216), .c(n323), .d(n172) );
	inv_2 U168 ( .x(n178), .a(n324) );
	exnor2_1 U169 ( .x(SUM[5]), .a(n178), .b(n103) );
	exnor2_1 U170 ( .x(SUM[19]), .a(n127), .b(n196) );
	exor2_1 U171 ( .x(SUM[4]), .a(n179), .b(n171) );
	exor2_1 U172 ( .x(n184), .a(A[28]), .b(B[28]) );
	exnor2_1 U173 ( .x(SUM[28]), .a(n183), .b(n184) );
	exnor2_1 U174 ( .x(SUM[8]), .a(n174), .b(n175) );
	inv_2 U175 ( .x(n230), .a(B[27]) );
	inv_2 U176 ( .x(n229), .a(A[27]) );
	inv_0 U177 ( .x(n63), .a(n364) );
	exnor2_1 U178 ( .x(SUM[9]), .a(n173), .b(n94) );
	exor2_1 U179 ( .x(SUM[15]), .a(n200), .b(n201) );
	inv_2 U18 ( .x(n306), .a(n151) );
	inv_2 U180 ( .x(n160), .a(n75) );
	exnor2_1 U181 ( .x(SUM[21]), .a(n160), .b(n193) );
	exor2_1 U182 ( .x(SUM[23]), .a(n191), .b(n192) );
	oai211_1 U183 ( .x(n191), .a(n75), .b(n300), .c(n348), .d(n347) );
	exor2_1 U184 ( .x(n192), .a(A[23]), .b(B[23]) );
	exnor2_1 U185 ( .x(SUM[24]), .a(n189), .b(n190) );
	exor2_1 U186 ( .x(n188), .a(B[25]), .b(A[25]) );
	exnor2_1 U187 ( .x(SUM[25]), .a(n93), .b(n188) );
	exnor2_1 U188 ( .x(SUM[29]), .a(n64), .b(n52) );
	inv_2 U189 ( .x(n209), .a(B[1]) );
	inv_2 U19 ( .x(n210), .a(n58) );
	nand4_2 U190 ( .x(n219), .a(n220), .b(n221), .c(n222), .d(n223) );
	ao21_3 U191 ( .x(n51), .a(n165), .b(n80), .c(n166) );
	nand2i_3 U192 ( .x(n279), .a(B[18]), .b(n260) );
	exnor2_1 U193 ( .x(n52), .a(B[29]), .b(A[29]) );
	nor2_1 U194 ( .x(n112), .a(A[17]), .b(B[17]) );
	oai21_1 U195 ( .x(n197), .a(n199), .b(n133), .c(n132) );
	ao21_3 U197 ( .x(n53), .a(n80), .b(n162), .c(n164) );
	nand2i_0 U198 ( .x(n162), .a(B[29]), .b(n227) );
	nand3i_1 U20 ( .x(n223), .a(n284), .b(n310), .c(n287) );
	ao21_4 U200 ( .x(n329), .a(n56), .b(n55), .c(n54) );
	inv_3 U201 ( .x(n55), .a(n219) );
	nand3_1 U202 ( .x(n56), .a(n150), .b(n315), .c(n306) );
	inv_4 U203 ( .x(n356), .a(n254) );
	and3i_4 U204 ( .x(n153), .a(n151), .b(n154), .c(n315) );
	nand3_5 U205 ( .x(n151), .a(n210), .b(n211), .c(n212) );
	nor2i_1 U206 ( .x(n146), .a(n147), .b(n148) );
	inv_2 U208 ( .x(n215), .a(B[6]) );
	nand2i_2 U209 ( .x(n244), .a(A[13]), .b(n264) );
	nand2_0 U21 ( .x(n98), .a(A[7]), .b(B[7]) );
	nand2i_2 U210 ( .x(n243), .a(B[14]), .b(n265) );
	nand2i_2 U211 ( .x(n363), .a(A[15]), .b(n263) );
	nor2_1 U213 ( .x(n157), .a(n111), .b(n135) );
	inv_1 U214 ( .x(n259), .a(A[17]) );
	nand2_0 U215 ( .x(n369), .a(B[1]), .b(A[1]) );
	nand2_0 U216 ( .x(n358), .a(B[1]), .b(A[1]) );
	inv_2 U217 ( .x(n208), .a(A[1]) );
	nand2_1 U218 ( .x(n362), .a(B[1]), .b(A[1]) );
	nor2_2 U219 ( .x(n149), .a(B[1]), .b(A[1]) );
	nand4_1 U22 ( .x(n221), .a(n287), .b(n310), .c(n316), .d(n285) );
	aoi21_3 U220 ( .x(n167), .a(n168), .b(n163), .c(n166) );
	nand2_1 U221 ( .x(n252), .a(n57), .b(n256) );
	inv_1 U222 ( .x(n256), .a(A[10]) );
	exnor2_1 U223 ( .x(SUM[20]), .a(n194), .b(n195) );
	nand2_0 U224 ( .x(n172), .a(B[4]), .b(A[4]) );
	inv_12 U225 ( .x(n216), .a(A[4]) );
	or2_2 U226 ( .x(n147), .a(n256), .b(n84) );
	inv_2 U227 ( .x(n214), .a(B[5]) );
	nand2_5 U228 ( .x(n58), .a(n310), .b(n287) );
	nand2i_2 U23 ( .x(n316), .a(A[5]), .b(n214) );
	inv_1 U230 ( .x(n257), .a(A[11]) );
	exor2_1 U231 ( .x(n201), .a(A[15]), .b(B[15]) );
	aoi21_1 U232 ( .x(n276), .a(A[15]), .b(B[15]), .c(n157) );
	nand4_3 U233 ( .x(n336), .a(n339), .b(n338), .c(n337), .d(n340) );
	inv_0 U234 ( .x(n59), .a(n278) );
	inv_2 U235 ( .x(n60), .a(n59) );
	nand2_0 U236 ( .x(n289), .a(A[8]), .b(B[8]) );
	inv_0 U237 ( .x(n225), .a(A[8]) );
	inv_7 U238 ( .x(n213), .a(A[7]) );
	oai211_3 U239 ( .x(n339), .a(n219), .b(n153), .c(n357), .d(n356) );
	inv_10 U240 ( .x(n357), .a(n247) );
	inv_2 U242 ( .x(n194), .a(n336) );
	nor2i_0 U243 ( .x(n128), .a(n279), .b(n239) );
	oaoi211_2 U244 ( .x(n76), .a(n79), .b(n78), .c(n336), .d(n77) );
	aoai211_1 U245 ( .x(n189), .a(n267), .b(n266), .c(n75), .d(n353) );
	inv_2 U246 ( .x(n62), .a(n180) );
	exor2_1 U247 ( .x(n180), .a(B[31]), .b(A[31]) );
	aoai211_1 U248 ( .x(n64), .a(n268), .b(n269), .c(n63), .d(n346) );
	nand4i_1 U249 ( .x(n220), .a(n152), .b(n310), .c(n287), .d(n286) );
	nor2_1 U25 ( .x(n286), .a(n170), .b(n118) );
	nand2_1 U250 ( .x(n308), .a(B[17]), .b(A[17]) );
	exor2_1 U251 ( .x(SUM[27]), .a(n82), .b(n186) );
	ao221_4 U252 ( .x(n80), .a(n364), .b(n87), .c(n364), .d(n86), .e(n85) );
	inv_0 U253 ( .x(n65), .a(n255) );
	nand2i_2 U254 ( .x(n352), .a(n95), .b(n89) );
	nand3i_1 U255 ( .x(n326), .a(n289), .b(n251), .c(n89) );
	inv_0 U256 ( .x(n148), .a(n89) );
	nand2_1 U257 ( .x(n309), .a(A[16]), .b(B[16]) );
	mx4_4 U258 ( .x(n185), .d0(B[26]), .sl0(A[26]), .d1(n361), .sl1(n66), .d2(n344),
		.sl2(n67), .d3(n361), .sl3(n68) );
	inv_2 U259 ( .x(n66), .a(n298) );
	inv_2 U260 ( .x(n67), .a(n116) );
	inv_2 U261 ( .x(n68), .a(n297) );
	oaoi211_1 U262 ( .x(n71), .a(n69), .b(n260), .c(n278), .d(n70) );
	inv_7 U263 ( .x(n260), .a(A[18]) );
	nand2_4 U264 ( .x(n125), .a(B[2]), .b(A[2]) );
	ao21_2 U265 ( .x(n278), .a(n308), .b(n309), .c(n112) );
	nand2i_6 U266 ( .x(n315), .a(B[2]), .b(n207) );
	nand2_0 U268 ( .x(n104), .a(B[5]), .b(A[5]) );
	nand2_0 U269 ( .x(n284), .a(B[5]), .b(A[5]) );
	inv_2 U27 ( .x(n54), .a(n356) );
	nor2_0 U270 ( .x(n152), .a(A[5]), .b(B[5]) );
	inv_2 U271 ( .x(n72), .a(n270) );
	inv_2 U272 ( .x(n73), .a(n271) );
	inv_0 U273 ( .x(n270), .a(B[30]) );
	inv_2 U274 ( .x(n271), .a(A[30]) );
	nand2_2 U275 ( .x(n305), .a(n306), .b(n307) );
	buf_3 U276 ( .x(n74), .a(n215) );
	inv_2 U279 ( .x(n77), .a(n350) );
	aoi21_1 U28 ( .x(n302), .a(n301), .b(n303), .c(n304) );
	inv_2 U280 ( .x(n78), .a(n237) );
	inv_2 U281 ( .x(n79), .a(n236) );
	nand2_0 U282 ( .x(n350), .a(A[20]), .b(B[20]) );
	inv_0 U283 ( .x(n237), .a(A[20]) );
	inv_0 U284 ( .x(n236), .a(B[20]) );
	nor2_0 U285 ( .x(n156), .a(B[1]), .b(A[1]) );
	nor2i_0 U286 ( .x(n124), .a(n125), .b(n126) );
	inv_2 U287 ( .x(n317), .a(n125) );
	oai211_1 U288 ( .x(n150), .a(n156), .b(n123), .c(n125), .d(n358) );
	aoai211_5 U289 ( .x(n364), .a(n229), .b(n230), .c(n345), .d(n351) );
	nor2_0 U29 ( .x(n301), .a(n142), .b(n145) );
	nand2_0 U290 ( .x(n343), .a(A[24]), .b(B[24]) );
	exor2_1 U291 ( .x(n198), .a(B[17]), .b(A[17]) );
	inv_0 U292 ( .x(n327), .a(n219) );
	ao21_1 U293 ( .x(n175), .a(A[8]), .b(B[8]), .c(n250) );
	inv_0 U294 ( .x(n82), .a(n345) );
	inv_3 U295 ( .x(n226), .a(B[9]) );
	nand2_2 U296 ( .x(n95), .a(B[9]), .b(A[9]) );
	ao221_4 U297 ( .x(n163), .a(n364), .b(n87), .c(n364), .d(n86), .e(n85) );
	nor2_0 U298 ( .x(n169), .a(A[4]), .b(B[4]) );
	aoai211_1 U299 ( .x(n83), .a(n360), .b(n359), .c(n75), .d(n294) );
	inv_0 U30 ( .x(n145), .a(n253) );
	inv_0 U300 ( .x(n84), .a(B[10]) );
	inv_2 U301 ( .x(n85), .a(n346) );
	inv_2 U302 ( .x(n86), .a(n269) );
	inv_2 U303 ( .x(n87), .a(n268) );
	inv_0 U304 ( .x(n183), .a(n364) );
	nand2_0 U305 ( .x(n346), .a(B[28]), .b(A[28]) );
	inv_0 U306 ( .x(n269), .a(B[28]) );
	inv_0 U307 ( .x(n268), .a(A[28]) );
	nand2_2 U308 ( .x(n109), .a(B[21]), .b(A[21]) );
	nand2_0 U309 ( .x(n132), .a(A[16]), .b(B[16]) );
	inv_0 U31 ( .x(n264), .a(B[13]) );
	and2_2 U310 ( .x(n88), .a(A[6]), .b(B[6]) );
	inv_0 U311 ( .x(n101), .a(n88) );
	nand2_1 U312 ( .x(n138), .a(B[13]), .b(A[13]) );
	inv_4 U313 ( .x(n238), .a(B[12]) );
	nor3i_5 U314 ( .x(n115), .a(n116), .b(n92), .c(n114) );
	exnor2_5 U315 ( .x(SUM[26]), .a(n115), .b(n187) );
	inv_6 U316 ( .x(n207), .a(A[2]) );
	nand2i_4 U317 ( .x(n245), .a(n70), .b(n374) );
	or3i_5 U318 ( .x(n247), .a(n248), .b(n113), .c(n241) );
	nand2i_4 U319 ( .x(n254), .a(n142), .b(n255) );
	nand2_3 U32 ( .x(n203), .a(n302), .b(n329) );
	inv_6 U320 ( .x(n265), .a(A[14]) );
	oai21_4 U321 ( .x(n274), .a(n242), .b(n275), .c(n276) );
	exnor2_3 U322 ( .x(n280), .a(n281), .b(n260) );
	mux2i_3 U323 ( .x(SUM[22]), .d0(n120), .sl(n158), .d1(n282) );
	nor2i_5 U324 ( .x(n285), .a(B[4]), .b(n216) );
	nand2_2 U325 ( .x(n290), .a(n144), .b(n147) );
	oai21_4 U326 ( .x(n292), .a(n261), .b(n262), .c(n293) );
	nand2_2 U327 ( .x(n164), .a(n299), .b(n271) );
	exor2_3 U328 ( .x(n181), .a(B[30]), .b(n73) );
	exor2_3 U329 ( .x(n187), .a(A[26]), .b(B[26]) );
	nand2_1 U33 ( .x(n331), .a(n203), .b(n244) );
	nand2i_4 U330 ( .x(n211), .a(B[3]), .b(n218) );
	nand3i_3 U331 ( .x(n307), .a(n317), .b(n320), .c(n319) );
	inv_5 U334 ( .x(n345), .a(n185) );
	oai21_4 U335 ( .x(n206), .a(n173), .b(n96), .c(n95) );
	inv_5 U336 ( .x(n349), .a(n206) );
	nand2i_4 U337 ( .x(n340), .a(n141), .b(n357) );
	nand3i_3 U338 ( .x(n338), .a(n291), .b(n303), .c(n357) );
	nand2i_4 U339 ( .x(n359), .a(n342), .b(n355) );
	nand3_1 U34 ( .x(n241), .a(n363), .b(n243), .c(n244) );
	aoai211_4 U340 ( .x(n337), .a(n248), .b(n274), .c(n292), .d(n335) );
	mux2i_3 U341 ( .x(n90), .d0(n283), .sl(B[18]), .d1(n280) );
	nand2_3 U342 ( .x(SUM[18]), .a(n90), .b(n91) );
	nand2i_6 U344 ( .x(n159), .a(A[21]), .b(n233) );
	nor2i_5 U345 ( .x(n92), .a(B[25]), .b(n93) );
	nor2i_5 U346 ( .x(n114), .a(A[25]), .b(n93) );
	nand2i_6 U347 ( .x(n251), .a(A[9]), .b(n226) );
	nand2i_5 U348 ( .x(n333), .a(n241), .b(n203) );
	inv_10 U349 ( .x(n217), .a(B[4]) );
	inv_2 U35 ( .x(n258), .a(A[16]) );
	nand2i_6 U350 ( .x(n310), .a(A[6]), .b(n74) );
	nand2i_6 U351 ( .x(n287), .a(B[7]), .b(n213) );
	aoi21_4 U352 ( .x(n222), .a(n88), .b(n287), .c(n288) );
	inv_6 U353 ( .x(n248), .a(n245) );
	nand2i_4 U354 ( .x(n291), .a(n142), .b(n253) );
	aoi21_4 U355 ( .x(n212), .a(n217), .b(n216), .c(n105) );
	inv_16 U356 ( .x(n262), .a(A[19]) );
	nor2_8 U357 ( .x(n113), .a(A[19]), .b(B[19]) );
	nor2i_1 U358 ( .x(n283), .a(A[18]), .b(n277) );
	oai21_3 U359 ( .x(n277), .a(n199), .b(n239), .c(n60) );
	nand2_2 U36 ( .x(n273), .a(A[23]), .b(B[23]) );
	inv_0 U360 ( .x(n370), .a(n105) );
	inv_2 U361 ( .x(n371), .a(n370) );
	inv_3 U362 ( .x(n105), .a(n316) );
	exnor2_1 U363 ( .x(SUM[11]), .a(n205), .b(n372) );
	inv_2 U364 ( .x(n372), .a(n143) );
	oai21_2 U365 ( .x(n205), .a(n148), .b(n349), .c(n147) );
	nor2i_0 U366 ( .x(n143), .a(n144), .b(n373) );
	oai211_1 U367 ( .x(n154), .a(n149), .b(n123), .c(n125), .d(n362) );
	nand2_3 U368 ( .x(n123), .a(B[0]), .b(A[0]) );
	oaoi211_2 U369 ( .x(n75), .a(n79), .b(n78), .c(n61), .d(n77) );
	nor2_1 U37 ( .x(n110), .a(A[23]), .b(B[23]) );
	inv_4 U370 ( .x(n61), .a(n194) );
	nand2_1 U371 ( .x(n174), .a(n81), .b(n305) );
	inv_2 U372 ( .x(n81), .a(n219) );
	inv_0 U373 ( .x(n373), .a(n253) );
	nand2i_3 U374 ( .x(n253), .a(B[11]), .b(n257) );
	inv_4 U375 ( .x(n255), .a(n249) );
	nand4i_3 U376 ( .x(n249), .a(n250), .b(n251), .c(n89), .d(n253) );
	buf_6 U377 ( .x(n89), .a(n252) );
	nor2i_3 U378 ( .x(n374), .a(n334), .b(n375) );
	inv_0 U379 ( .x(n239), .a(n374) );
	nor2i_1 U38 ( .x(n108), .a(n109), .b(n106) );
	inv_5 U380 ( .x(n375), .a(n240) );
	inv_0 U381 ( .x(n133), .a(n334) );
	nand2i_2 U382 ( .x(n240), .a(B[17]), .b(n259) );
	nand2i_2 U383 ( .x(n334), .a(B[16]), .b(n258) );
	aoai211_3 U384 ( .x(n361), .a(n360), .b(n359), .c(n76), .d(n294) );
	nor2i_1 U39 ( .x(n106), .a(A[22]), .b(n107) );
	inv_2 U40 ( .x(n107), .a(B[22]) );
	nand3i_1 U41 ( .x(n319), .a(n149), .b(n315), .c(n318) );
	or3i_2 U42 ( .x(n320), .a(n315), .b(n209), .c(n208) );
	inv_2 U43 ( .x(n126), .a(n315) );
	aoi21_1 U44 ( .x(n122), .a(n123), .b(n369), .c(n367) );
	nand2i_2 U45 ( .x(n313), .a(B[1]), .b(n208) );
	inv_2 U46 ( .x(n318), .a(n123) );
	nand2i_2 U47 ( .x(n312), .a(A[12]), .b(n238) );
	inv_2 U48 ( .x(n142), .a(n312) );
	nand2_0 U49 ( .x(n141), .a(A[12]), .b(B[12]) );
	exnor2_3 U5 ( .x(SUM[31]), .a(n50), .b(n49) );
	nor2i_1 U50 ( .x(n140), .a(n141), .b(n142) );
	nand2i_2 U51 ( .x(n328), .a(n373), .b(n303) );
	aoai211_1 U53 ( .x(n204), .a(n327), .b(n305), .c(n65), .d(n328) );
	inv_2 U54 ( .x(n288), .a(n98) );
	nand2i_2 U55 ( .x(n297), .a(n155), .b(B[25]) );
	nand2i_2 U56 ( .x(n298), .a(n155), .b(A[25]) );
	nand2i_2 U57 ( .x(n344), .a(B[26]), .b(n231) );
	inv_2 U58 ( .x(n231), .a(A[26]) );
	inv_2 U59 ( .x(n155), .a(n344) );
	inv_2 U6 ( .x(n49), .a(n62) );
	nor2i_1 U60 ( .x(SUM[0]), .a(n365), .b(n366) );
	nor2_1 U61 ( .x(n366), .a(B[0]), .b(A[0]) );
	nand2_1 U62 ( .x(n144), .a(A[11]), .b(B[11]) );
	inv_2 U64 ( .x(n304), .a(n141) );
	nand2i_2 U65 ( .x(n335), .a(B[19]), .b(n262) );
	inv_2 U66 ( .x(n261), .a(B[19]) );
	nand3i_2 U67 ( .x(n303), .a(n290), .b(n352), .c(n326) );
	nand2_1 U68 ( .x(n135), .a(A[14]), .b(B[14]) );
	nor2i_1 U69 ( .x(n134), .a(n135), .b(n136) );
	aoi22_1 U7 ( .x(n50), .a(n51), .b(n73), .c(n53), .d(n72) );
	exor2_1 U70 ( .x(SUM[13]), .a(n203), .b(n137) );
	nor2i_1 U71 ( .x(n137), .a(n138), .b(n139) );
	inv_2 U72 ( .x(n139), .a(n244) );
	inv_1 U73 ( .x(n57), .a(B[10]) );
	aoi21_1 U74 ( .x(n158), .a(n159), .b(n160), .c(n161) );
	exnor2_1 U75 ( .x(n282), .a(A[22]), .b(B[22]) );
	aoi21_1 U76 ( .x(n120), .a(A[22]), .b(B[22]), .c(n121) );
	inv_3 U77 ( .x(n121), .a(n314) );
	exor2_1 U78 ( .x(n196), .a(A[19]), .b(B[19]) );
	inv_2 U79 ( .x(n70), .a(n279) );
	nand2i_2 U8 ( .x(n311), .a(A[8]), .b(n224) );
	inv_0 U80 ( .x(n69), .a(B[18]) );
	inv_2 U81 ( .x(n293), .a(n71) );
	inv_0 U82 ( .x(n130), .a(n293) );
	nand2i_3 U83 ( .x(n129), .a(n274), .b(n333) );
	aoi21_1 U84 ( .x(n127), .a(n128), .b(n129), .c(n130) );
	nor2i_1 U85 ( .x(n171), .a(n172), .b(n169) );
	oai21_1 U86 ( .x(n179), .a(n119), .b(n182), .c(n118) );
	inv_0 U87 ( .x(n218), .a(A[3]) );
	nand2_1 U88 ( .x(n118), .a(A[3]), .b(B[3]) );
	nand2i_0 U89 ( .x(n91), .a(n279), .b(n277) );
	inv_3 U9 ( .x(n224), .a(B[8]) );
	inv_2 U90 ( .x(n281), .a(n277) );
	inv_2 U91 ( .x(n228), .a(B[29]) );
	nand2i_2 U92 ( .x(n168), .a(A[29]), .b(n228) );
	nand2_2 U93 ( .x(n351), .a(B[27]), .b(A[27]) );
	nand2i_2 U94 ( .x(n165), .a(B[29]), .b(n227) );
	inv_2 U95 ( .x(n227), .a(A[29]) );
	inv_2 U96 ( .x(n166), .a(n299) );
	nand2_2 U97 ( .x(n299), .a(B[29]), .b(A[29]) );
	exnor2_1 U98 ( .x(SUM[1]), .a(n368), .b(n365) );
	nor2i_1 U99 ( .x(n368), .a(n369), .b(n367) );

endmodule


module EX_DW01_add_32_6_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
	n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
	n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
	n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
	n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
	n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
	n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
	n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
	n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
	n352, n353, n354, n355, n356, n357, n358, n359, n361, n362, n363, n364,
	n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
	n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n49, n50,
	n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
	n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
	n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
	n93, n94, n95, n96, n97, n98, n99;


	ao211_2 U10 ( .x(n350), .a(n89), .b(n239), .c(n241), .d(n240) );
	inv_2 U100 ( .x(n336), .a(n147) );
	nand2_1 U101 ( .x(n147), .a(B[2]), .b(A[2]) );
	nand3_3 U102 ( .x(n367), .a(n84), .b(n366), .c(n54) );
	inv_2 U103 ( .x(n140), .a(B[26]) );
	nor2i_1 U104 ( .x(n139), .a(A[26]), .b(n140) );
	nand2i_2 U105 ( .x(n200), .a(n56), .b(n255) );
	nand2_2 U106 ( .x(n331), .a(n56), .b(A[29]) );
	inv_2 U107 ( .x(n255), .a(A[29]) );
	nand2i_2 U108 ( .x(n204), .a(n56), .b(n255) );
	oai21_1 U109 ( .x(n298), .a(A[1]), .b(B[1]), .c(n342) );
	inv_0 U11 ( .x(n190), .a(n350) );
	exor2_1 U110 ( .x(SUM[1]), .a(n298), .b(n384) );
	nor2i_1 U111 ( .x(n153), .a(n154), .b(n155) );
	inv_2 U112 ( .x(n79), .a(n275) );
	inv_2 U113 ( .x(n155), .a(n361) );
	inv_0 U114 ( .x(n260), .a(B[21]) );
	inv_2 U115 ( .x(n363), .a(n196) );
	nand2i_2 U116 ( .x(n227), .a(n363), .b(n132) );
	exor2_1 U117 ( .x(n226), .a(A[23]), .b(B[23]) );
	oai211_1 U118 ( .x(n225), .a(n82), .b(n278), .c(n371), .d(n370) );
	nand2i_2 U119 ( .x(n370), .a(n145), .b(n198) );
	buf_1 U12 ( .x(n50), .a(n164) );
	inv_2 U120 ( .x(n198), .a(n132) );
	exnor2_1 U121 ( .x(SUM[24]), .a(n223), .b(n224) );
	inv_0 U122 ( .x(n379), .a(n288) );
	nand2i_2 U123 ( .x(n224), .a(n364), .b(n365) );
	inv_2 U124 ( .x(n364), .a(n326) );
	exor2_1 U125 ( .x(n222), .a(n54), .b(A[25]) );
	exor2_1 U126 ( .x(n220), .a(A[26]), .b(B[26]) );
	nand2_2 U127 ( .x(n188), .a(A[25]), .b(n54) );
	inv_2 U128 ( .x(n283), .a(A[25]) );
	inv_2 U129 ( .x(n282), .a(n54) );
	nand2_0 U13 ( .x(n289), .a(A[23]), .b(B[23]) );
	exnor2_1 U130 ( .x(SUM[3]), .a(n51), .b(n141) );
	exor2_1 U131 ( .x(SUM[2]), .a(n230), .b(n146) );
	oai21_1 U132 ( .x(n230), .a(n384), .b(n181), .c(n342) );
	inv_7 U133 ( .x(n181), .a(n382) );
	nor2i_1 U134 ( .x(n146), .a(n147), .b(n148) );
	inv_2 U135 ( .x(n148), .a(n302) );
	exor2_1 U136 ( .x(SUM[12]), .a(n236), .b(n166) );
	nor2i_1 U138 ( .x(n166), .a(n167), .b(n168) );
	nor2i_1 U14 ( .x(n131), .a(n132), .b(n129) );
	exnor2_1 U140 ( .x(SUM[7]), .a(n115), .b(n118) );
	exor2_1 U141 ( .x(SUM[11]), .a(n237), .b(n169) );
	ao21_2 U142 ( .x(n237), .a(n238), .b(n103), .c(n344) );
	nor2i_1 U143 ( .x(n169), .a(n170), .b(n171) );
	exor2_1 U144 ( .x(n229), .a(A[20]), .b(B[20]) );
	exor2_1 U145 ( .x(SUM[14]), .a(n157), .b(n160) );
	oai21_1 U146 ( .x(n157), .a(n165), .b(n372), .c(n50) );
	nor2i_1 U147 ( .x(n160), .a(n161), .b(n162) );
	inv_0 U148 ( .x(n162), .a(n158) );
	inv_2 U149 ( .x(n372), .a(n235) );
	nand2i_2 U15 ( .x(n378), .a(n318), .b(n307) );
	nor2i_1 U150 ( .x(n163), .a(n50), .b(n165) );
	inv_2 U151 ( .x(n168), .a(n275) );
	oai21_1 U152 ( .x(n235), .a(n386), .b(n168), .c(n167) );
	exor2_1 U153 ( .x(SUM[13]), .a(n235), .b(n163) );
	exor2_1 U154 ( .x(SUM[10]), .a(n238), .b(n172) );
	mux2i_1 U155 ( .x(SUM[22]), .d0(n144), .sl(n195), .d1(n299) );
	exor2_1 U156 ( .x(SUM[5]), .a(n211), .b(n123) );
	aoi21_1 U157 ( .x(n85), .a(n348), .b(n212), .c(n86) );
	nor2i_1 U158 ( .x(n123), .a(n124), .b(n125) );
	exnor2_1 U159 ( .x(SUM[19]), .a(n149), .b(n231) );
	inv_6 U16 ( .x(n107), .a(A[6]) );
	exor2_1 U160 ( .x(SUM[4]), .a(n212), .b(n126) );
	oai21_1 U161 ( .x(n212), .a(n143), .b(n51), .c(n142) );
	nand2_2 U162 ( .x(SUM[18]), .a(n110), .b(n111) );
	mux2i_1 U163 ( .x(n110), .d0(n300), .sl(B[18]), .d1(n296) );
	nand2i_2 U164 ( .x(n111), .a(n295), .b(n292) );
	exnor2_3 U165 ( .x(SUM[30]), .a(n206), .b(n214) );
	exor2_1 U166 ( .x(n216), .a(A[28]), .b(B[28]) );
	exnor2_1 U167 ( .x(SUM[8]), .a(n209), .b(n210) );
	oai211_1 U168 ( .x(n209), .a(n51), .b(n61), .c(n351), .d(n305) );
	exor2_1 U169 ( .x(n215), .a(n56), .b(A[29]) );
	inv_0 U17 ( .x(n62), .a(B[2]) );
	inv_2 U170 ( .x(n286), .a(B[30]) );
	inv_2 U171 ( .x(n287), .a(A[30]) );
	exnor2_1 U172 ( .x(SUM[9]), .a(n208), .b(n112) );
	oai22_1 U173 ( .x(n353), .a(n252), .b(n253), .c(n313), .d(n352) );
	inv_5 U174 ( .x(n313), .a(n346) );
	inv_2 U175 ( .x(n352), .a(n209) );
	nor2i_0 U176 ( .x(n112), .a(n113), .b(n114) );
	inv_2 U177 ( .x(n159), .a(n161) );
	aoi21_1 U178 ( .x(n156), .a(n157), .b(n158), .c(n159) );
	exnor2_1 U179 ( .x(SUM[15]), .a(n156), .b(n234) );
	aoai211_1 U18 ( .x(n100), .a(n99), .b(n265), .c(n164), .d(n310) );
	exnor2_1 U180 ( .x(SUM[16]), .a(n77), .b(n153) );
	exor2_1 U181 ( .x(SUM[23]), .a(n225), .b(n226) );
	exnor2_1 U182 ( .x(SUM[25]), .a(n221), .b(n222) );
	exor2_1 U183 ( .x(SUM[29]), .a(n201), .b(n215) );
	oa211_2 U184 ( .x(n51), .a(n384), .b(n301), .c(n350), .d(n147) );
	exnor2_1 U186 ( .x(n52), .a(B[31]), .b(A[31]) );
	inv_2 U187 ( .x(n143), .a(n347) );
	nand2i_2 U188 ( .x(n347), .a(B[3]), .b(n249) );
	inv_2 U189 ( .x(n128), .a(n348) );
	inv_5 U19 ( .x(n315), .a(n312) );
	nand2_2 U190 ( .x(n348), .a(n93), .b(n246) );
	buf_3 U191 ( .x(n54), .a(B[25]) );
	inv_0 U192 ( .x(n55), .a(B[29]) );
	inv_2 U193 ( .x(n56), .a(n55) );
	inv_2 U194 ( .x(n58), .a(n81) );
	inv_6 U195 ( .x(n245), .a(A[5]) );
	aoi21_2 U196 ( .x(n57), .a(n228), .b(n83), .c(n106) );
	aoai211_3 U197 ( .x(n84), .a(n381), .b(n380), .c(n57), .d(n325) );
	aoi21_2 U198 ( .x(n325), .a(n288), .b(n326), .c(n327) );
	and3i_1 U20 ( .x(n192), .a(n174), .b(A[9]), .c(B[9]) );
	inv_2 U200 ( .x(n106), .a(n373) );
	nand2_4 U201 ( .x(n60), .a(n59), .b(n262) );
	inv_4 U202 ( .x(n59), .a(B[17]) );
	inv_7 U203 ( .x(n262), .a(A[17]) );
	inv_5 U204 ( .x(n261), .a(A[16]) );
	inv_1 U205 ( .x(n75), .a(B[10]) );
	nand2_2 U207 ( .x(n142), .a(A[3]), .b(B[3]) );
	nand3_1 U208 ( .x(n61), .a(n243), .b(n244), .c(n347) );
	nor2_3 U209 ( .x(n243), .a(n53), .b(n120) );
	nor2i_0 U21 ( .x(n134), .a(B[18]), .b(n135) );
	nand3_2 U210 ( .x(n242), .a(n243), .b(n244), .c(n347) );
	nand2i_3 U211 ( .x(n349), .a(B[5]), .b(n245) );
	oa22_4 U212 ( .x(n77), .a(n273), .b(n175), .c(n386), .d(n185) );
	nand2i_3 U213 ( .x(n355), .a(A[15]), .b(n268) );
	and4i_4 U214 ( .x(n78), .a(n79), .b(n355), .c(n274), .d(n158) );
	inv_2 U215 ( .x(n273), .a(n355) );
	ao21_6 U216 ( .x(n314), .a(n62), .b(n239), .c(n315) );
	aoai211_3 U217 ( .x(n201), .a(n284), .b(n285), .c(n63), .d(n369) );
	nand3i_5 U218 ( .x(n217), .a(n139), .b(n367), .c(n329) );
	aoai211_3 U219 ( .x(n64), .a(n381), .b(n380), .c(n105), .d(n325) );
	inv_8 U22 ( .x(n135), .a(A[18]) );
	aoai211_1 U220 ( .x(n330), .a(n381), .b(n380), .c(n58), .d(n325) );
	and3i_3 U221 ( .x(n183), .a(n193), .b(n66), .c(n65) );
	inv_2 U222 ( .x(n65), .a(n192) );
	or3_5 U223 ( .x(n66), .a(n174), .b(n114), .c(n194) );
	nand2_2 U224 ( .x(n193), .a(n170), .b(n173) );
	inv_2 U225 ( .x(n279), .a(n67) );
	inv_2 U226 ( .x(n68), .a(B[23]) );
	inv_0 U227 ( .x(n280), .a(n278) );
	ao31_6 U228 ( .x(n95), .a(n176), .b(n161), .c(n177), .d(n178) );
	nor2i_3 U229 ( .x(n319), .a(A[4]), .b(n320) );
	inv_5 U23 ( .x(n97), .a(B[16]) );
	inv_5 U230 ( .x(n93), .a(A[4]) );
	buf_1 U231 ( .x(n69), .a(n228) );
	nand2i_2 U233 ( .x(n306), .a(B[5]), .b(n245) );
	ao21_4 U234 ( .x(n238), .a(n353), .b(n71), .c(n70) );
	inv_2 U235 ( .x(n70), .a(n113) );
	inv_0 U236 ( .x(n71), .a(n114) );
	inv_0 U237 ( .x(n208), .a(n353) );
	aoi21_3 U238 ( .x(n329), .a(n64), .b(n328), .c(n186) );
	inv_5 U239 ( .x(n268), .a(B[15]) );
	nand2i_0 U24 ( .x(n290), .a(n270), .b(n291) );
	exor2_1 U240 ( .x(n234), .a(A[15]), .b(B[15]) );
	nand2_0 U241 ( .x(n339), .a(A[15]), .b(B[15]) );
	nand2_1 U242 ( .x(n310), .a(A[15]), .b(B[15]) );
	nor3_5 U243 ( .x(n316), .a(n189), .b(n314), .c(n242) );
	nand2_1 U244 ( .x(n119), .a(A[7]), .b(B[7]) );
	exor2_1 U245 ( .x(SUM[6]), .a(n116), .b(n121) );
	inv_0 U246 ( .x(n72), .a(n130) );
	or2_2 U247 ( .x(n365), .a(n73), .b(n74) );
	inv_1 U248 ( .x(n74), .a(B[24]) );
	and2_2 U249 ( .x(n179), .a(n75), .b(n76) );
	inv_3 U25 ( .x(n270), .a(n60) );
	inv_4 U250 ( .x(n241), .a(B[1]) );
	oai22_2 U251 ( .x(n213), .a(n203), .b(n287), .c(n199), .d(n286) );
	inv_6 U252 ( .x(n185), .a(n78) );
	and3_1 U253 ( .x(n175), .a(n80), .b(n176), .c(n375) );
	and2_1 U254 ( .x(n80), .a(n339), .b(n161) );
	nand2i_2 U255 ( .x(n275), .a(B[12]), .b(n266) );
	inv_1 U256 ( .x(n98), .a(B[17]) );
	inv_2 U257 ( .x(n82), .a(n81) );
	inv_2 U258 ( .x(n83), .a(n138) );
	nand4i_1 U259 ( .x(n381), .a(n145), .b(n196), .c(A[23]), .d(n326) );
	nand2_2 U26 ( .x(n291), .a(n97), .b(n261) );
	inv_14 U260 ( .x(n99), .a(B[14]) );
	exor2_1 U261 ( .x(SUM[20]), .a(n69), .b(n229) );
	nand3_4 U262 ( .x(n176), .a(n274), .b(n158), .c(n356) );
	nand2i_0 U263 ( .x(n375), .a(n164), .b(n158) );
	nand2i_4 U264 ( .x(n161), .a(n265), .b(B[14]) );
	aoai211_5 U265 ( .x(n383), .a(n256), .b(n257), .c(n368), .d(n374) );
	inv_10 U266 ( .x(n368), .a(n217) );
	inv_16 U267 ( .x(n265), .a(A[14]) );
	aoi31_1 U268 ( .x(n305), .a(n306), .b(n307), .c(n308), .d(n309) );
	nand4i_5 U269 ( .x(n324), .a(n309), .b(n351), .c(n377), .d(n378) );
	inv_2 U27 ( .x(n271), .a(n291) );
	inv_6 U270 ( .x(n309), .a(n376) );
	inv_0 U271 ( .x(n211), .a(n85) );
	inv_2 U272 ( .x(n86), .a(n127) );
	nand2_0 U273 ( .x(n127), .a(n109), .b(A[4]) );
	exor2_1 U274 ( .x(SUM[27]), .a(n217), .b(n218) );
	aoai211_2 U275 ( .x(n88), .a(n256), .b(n257), .c(n368), .d(n374) );
	inv_10 U276 ( .x(n240), .a(A[1]) );
	ao23_6 U277 ( .x(n362), .a(n137), .b(n264), .c(n95), .d(n340), .e(n94) );
	inv_2 U278 ( .x(n94), .a(n136) );
	inv_0 U279 ( .x(n264), .a(A[19]) );
	nor2_1 U28 ( .x(n186), .a(n187), .b(n188) );
	inv_2 U280 ( .x(n90), .a(B[7]) );
	inv_6 U281 ( .x(n250), .a(B[6]) );
	aoi21_3 U282 ( .x(n203), .a(n204), .b(n104), .c(n205) );
	inv_2 U283 ( .x(n205), .a(n331) );
	inv_0 U284 ( .x(n281), .a(n91) );
	nand2i_2 U286 ( .x(n178), .a(n273), .b(n311) );
	nand2i_6 U287 ( .x(n302), .a(B[2]), .b(n239) );
	aoai211_1 U288 ( .x(n223), .a(n281), .b(n279), .c(n82), .d(n379) );
	nand2i_2 U289 ( .x(n357), .a(B[10]), .b(n76) );
	nand2i_2 U29 ( .x(n366), .a(B[26]), .b(n258) );
	nor2i_0 U290 ( .x(n136), .a(A[19]), .b(n137) );
	nand2_0 U291 ( .x(n124), .a(B[5]), .b(A[5]) );
	nand2_0 U292 ( .x(n318), .a(B[5]), .b(A[5]) );
	aoi211_1 U293 ( .x(n96), .a(n262), .b(n98), .c(n261), .d(n97) );
	inv_0 U294 ( .x(n294), .a(n96) );
	nand2_1 U295 ( .x(n293), .a(B[17]), .b(A[17]) );
	nor2_5 U296 ( .x(n189), .a(n49), .b(n191) );
	inv_3 U297 ( .x(n177), .a(n100) );
	nor2i_0 U298 ( .x(n121), .a(n122), .b(n53) );
	nor2_2 U299 ( .x(n303), .a(n53), .b(n120) );
	inv_2 U30 ( .x(n258), .a(A[26]) );
	inv_0 U300 ( .x(n101), .a(n53) );
	nor2_0 U301 ( .x(n385), .a(B[0]), .b(A[0]) );
	inv_0 U302 ( .x(n102), .a(n357) );
	inv_2 U303 ( .x(n103), .a(n102) );
	oai21_3 U304 ( .x(n191), .a(n384), .b(n181), .c(n147) );
	nor2i_0 U305 ( .x(n126), .a(n127), .b(n128) );
	nand2i_2 U306 ( .x(n326), .a(B[24]), .b(n259) );
	exor2_1 U307 ( .x(n233), .a(B[17]), .b(A[17]) );
	ao221_4 U308 ( .x(n104), .a(n383), .b(A[28]), .c(n383), .d(B[28]), .e(n108) );
	nand2_2 U309 ( .x(n194), .a(A[8]), .b(B[8]) );
	inv_2 U31 ( .x(n187), .a(n366) );
	ao21_1 U310 ( .x(n210), .a(A[8]), .b(B[8]), .c(n313) );
	inv_0 U311 ( .x(n252), .a(B[8]) );
	nand2_0 U312 ( .x(n373), .a(A[20]), .b(B[20]) );
	nand2_0 U313 ( .x(n333), .a(A[9]), .b(B[9]) );
	inv_3 U314 ( .x(n254), .a(B[9]) );
	nand2_0 U315 ( .x(n113), .a(B[9]), .b(A[9]) );
	exnor2_1 U316 ( .x(SUM[28]), .a(n63), .b(n216) );
	aoi21_2 U317 ( .x(n199), .a(n200), .b(n104), .c(n202) );
	exnor2_3 U318 ( .x(SUM[31]), .a(n213), .b(n52) );
	inv_2 U319 ( .x(n108), .a(n369) );
	nand2_2 U32 ( .x(n374), .a(B[27]), .b(A[27]) );
	nand2_0 U320 ( .x(n369), .a(B[28]), .b(A[28]) );
	inv_0 U321 ( .x(n285), .a(B[28]) );
	inv_0 U322 ( .x(n284), .a(A[28]) );
	inv_0 U323 ( .x(n109), .a(n246) );
	nand2_2 U324 ( .x(n132), .a(B[21]), .b(A[21]) );
	nand2i_0 U325 ( .x(n361), .a(B[16]), .b(n261) );
	nand2_0 U326 ( .x(n154), .a(A[16]), .b(B[16]) );
	nor2i_0 U327 ( .x(n172), .a(n173), .b(n174) );
	oai211_1 U328 ( .x(n334), .a(n174), .b(n333), .c(n170), .d(n173) );
	inv_0 U329 ( .x(n344), .a(n173) );
	inv_0 U33 ( .x(n165), .a(n274) );
	nand2_2 U330 ( .x(n167), .a(A[12]), .b(B[12]) );
	nand2_0 U331 ( .x(n173), .a(A[10]), .b(B[10]) );
	nor3_4 U332 ( .x(n182), .a(n183), .b(n184), .c(n185) );
	exor2_3 U333 ( .x(SUM[26]), .a(n219), .b(n220) );
	exnor2_3 U334 ( .x(SUM[21]), .a(n197), .b(n227) );
	exor2_3 U335 ( .x(SUM[17]), .a(n232), .b(n233) );
	inv_6 U336 ( .x(n263), .a(B[18]) );
	inv_6 U337 ( .x(n266), .a(A[12]) );
	ao211_5 U338 ( .x(n269), .a(n135), .b(n263), .c(n270), .d(n271) );
	or3i_5 U339 ( .x(n276), .a(n277), .b(n179), .c(n114) );
	nand2_6 U34 ( .x(n158), .a(n99), .b(n265) );
	nand2i_4 U340 ( .x(n295), .a(B[18]), .b(n135) );
	exnor2_3 U341 ( .x(n296), .a(n297), .b(n135) );
	nand2i_4 U342 ( .x(n301), .a(n181), .b(n302) );
	nor2_5 U343 ( .x(n304), .a(n125), .b(n142) );
	nor2_5 U344 ( .x(n277), .a(n171), .b(n313) );
	nor3_4 U346 ( .x(n322), .a(n321), .b(n185), .c(n276) );
	aoi22_3 U347 ( .x(n323), .a(n316), .b(n317), .c(n324), .d(n322) );
	nand2_2 U348 ( .x(n202), .a(n331), .b(n287) );
	nand2i_4 U349 ( .x(n346), .a(B[8]), .b(n253) );
	nor2_0 U35 ( .x(n138), .a(A[20]), .b(B[20]) );
	oai221_3 U350 ( .x(n219), .a(n221), .b(n282), .c(n221), .d(n283), .e(n188) );
	nand2_2 U351 ( .x(n371), .a(A[22]), .b(n72) );
	oai21_4 U352 ( .x(n232), .a(n77), .b(n155), .c(n154) );
	nand2_8 U353 ( .x(n384), .a(A[0]), .b(B[0]) );
	nand3i_5 U354 ( .x(n228), .a(n182), .b(n362), .c(n323) );
	inv_6 U355 ( .x(n221), .a(n330) );
	inv_7 U356 ( .x(n174), .a(n357) );
	nand2i_6 U358 ( .x(n196), .a(A[21]), .b(n260) );
	nand3_4 U359 ( .x(n351), .a(n303), .b(n348), .c(n304) );
	nor2i_1 U36 ( .x(n91), .a(n280), .b(n92) );
	nand2i_6 U360 ( .x(n354), .a(A[9]), .b(n254) );
	nor2_6 U361 ( .x(n180), .a(n384), .b(n181) );
	nand2i_6 U363 ( .x(n345), .a(A[22]), .b(n130) );
	nor2i_5 U364 ( .x(n328), .a(A[25]), .b(n187) );
	inv_10 U365 ( .x(n256), .a(A[27]) );
	inv_8 U366 ( .x(n257), .a(B[27]) );
	inv_6 U367 ( .x(n307), .a(n247) );
	nand3_5 U368 ( .x(n377), .a(n307), .b(B[4]), .c(n319) );
	nand2i_6 U369 ( .x(n312), .a(A[19]), .b(n137) );
	nand2i_2 U37 ( .x(n278), .a(n145), .b(n196) );
	nor2_8 U371 ( .x(n133), .a(A[23]), .b(B[23]) );
	nand2i_6 U372 ( .x(n382), .a(B[1]), .b(n240) );
	nor2i_8 U373 ( .x(n129), .a(A[22]), .b(n130) );
	oa211_4 U374 ( .x(n386), .a(n335), .b(n337), .c(n358), .d(n359) );
	inv_0 U375 ( .x(n236), .a(n386) );
	nand2i_1 U376 ( .x(n337), .a(n276), .b(n338) );
	oai31_1 U377 ( .x(n335), .a(n190), .b(n336), .c(n180), .d(n302) );
	inv_5 U378 ( .x(n63), .a(n88) );
	aoi21_3 U379 ( .x(n206), .a(n207), .b(n201), .c(n205) );
	inv_2 U38 ( .x(n92), .a(A[23]) );
	nand3i_2 U380 ( .x(n184), .a(n171), .b(n312), .c(n311) );
	nand2i_2 U381 ( .x(n321), .a(n315), .b(n311) );
	and3i_4 U382 ( .x(n317), .a(n185), .b(n87), .c(n311) );
	inv_7 U383 ( .x(n311), .a(n269) );
	inv_4 U384 ( .x(n267), .a(B[13]) );
	aoi21_5 U385 ( .x(n105), .a(n228), .b(n83), .c(n106) );
	inv_2 U39 ( .x(n73), .a(A[24]) );
	inv_2 U40 ( .x(n327), .a(n365) );
	oai31_1 U41 ( .x(n288), .a(n131), .b(n145), .c(n133), .d(n289) );
	nand2_3 U42 ( .x(n380), .a(n67), .b(n326) );
	nor2_3 U43 ( .x(n67), .a(n278), .b(n68) );
	inv_5 U44 ( .x(n130), .a(B[22]) );
	inv_2 U45 ( .x(n259), .a(A[24]) );
	nor2i_1 U46 ( .x(n141), .a(n142), .b(n143) );
	nand2_0 U47 ( .x(n342), .a(B[1]), .b(A[1]) );
	or2_3 U48 ( .x(n122), .a(n107), .b(n250) );
	inv_4 U49 ( .x(n171), .a(n343) );
	nand2i_2 U5 ( .x(n248), .a(B[7]), .b(n251) );
	inv_5 U50 ( .x(n114), .a(n354) );
	nor2_0 U51 ( .x(n332), .a(n114), .b(n194) );
	aoai211_1 U52 ( .x(n359), .a(n332), .b(n103), .c(n334), .d(n343) );
	nand2i_2 U53 ( .x(n358), .a(n276), .b(n324) );
	inv_5 U54 ( .x(n239), .a(A[2]) );
	inv_1 U55 ( .x(n89), .a(B[2]) );
	nor2i_1 U57 ( .x(n118), .a(n119), .b(n120) );
	aoi21_1 U58 ( .x(n115), .a(n116), .b(n101), .c(n117) );
	oai21_1 U59 ( .x(n116), .a(n125), .b(n85), .c(n124) );
	ao22_3 U6 ( .x(n247), .a(n107), .b(n250), .c(n90), .d(n251) );
	inv_4 U60 ( .x(n125), .a(n349) );
	and2_3 U61 ( .x(n53), .a(n107), .b(n250) );
	inv_0 U62 ( .x(n117), .a(n122) );
	exor2_1 U63 ( .x(n218), .a(B[27]), .b(A[27]) );
	nor2i_1 U64 ( .x(SUM[0]), .a(n384), .b(n385) );
	inv_2 U65 ( .x(n272), .a(B[11]) );
	nand2i_3 U66 ( .x(n343), .a(A[11]), .b(n272) );
	nand2_0 U67 ( .x(n170), .a(A[11]), .b(B[11]) );
	inv_4 U68 ( .x(n87), .a(n276) );
	inv_2 U69 ( .x(n137), .a(B[19]) );
	inv_3 U7 ( .x(n251), .a(A[7]) );
	nand2i_3 U70 ( .x(n274), .a(A[13]), .b(n267) );
	nand2i_2 U71 ( .x(n164), .a(n267), .b(A[13]) );
	inv_2 U72 ( .x(n356), .a(n167) );
	inv_4 U73 ( .x(n253), .a(A[8]) );
	inv_2 U74 ( .x(n81), .a(n105) );
	inv_1 U75 ( .x(n197), .a(n58) );
	aoi21_1 U76 ( .x(n195), .a(n196), .b(n197), .c(n198) );
	exnor2_1 U77 ( .x(n299), .a(A[22]), .b(n72) );
	aoi21_1 U78 ( .x(n144), .a(A[22]), .b(n72), .c(n145) );
	inv_5 U79 ( .x(n145), .a(n345) );
	inv_4 U8 ( .x(n76), .a(A[10]) );
	exor2_1 U80 ( .x(n231), .a(A[19]), .b(B[19]) );
	aoi21_1 U81 ( .x(n149), .a(n150), .b(n151), .c(n152) );
	nor2i_1 U82 ( .x(n150), .a(n295), .b(n290) );
	inv_0 U83 ( .x(n151), .a(n77) );
	inv_0 U84 ( .x(n152), .a(n340) );
	oai31_1 U85 ( .x(n340), .a(n134), .b(n96), .c(n341), .d(n295) );
	inv_2 U86 ( .x(n341), .a(n293) );
	inv_2 U87 ( .x(n246), .a(B[4]) );
	nor2i_0 U88 ( .x(n300), .a(A[18]), .b(n292) );
	oai211_1 U89 ( .x(n292), .a(n77), .b(n290), .c(n293), .d(n294) );
	inv_2 U9 ( .x(n49), .a(n350) );
	inv_2 U90 ( .x(n297), .a(n292) );
	exor2_1 U91 ( .x(n214), .a(B[30]), .b(A[30]) );
	nand2i_2 U92 ( .x(n207), .a(A[29]), .b(n55) );
	inv_2 U93 ( .x(n320), .a(n306) );
	ao21_3 U94 ( .x(n376), .a(n119), .b(n122), .c(n120) );
	nand2_2 U95 ( .x(n308), .a(n127), .b(n124) );
	inv_5 U96 ( .x(n120), .a(n248) );
	aoi21_2 U97 ( .x(n244), .a(n93), .b(n246), .c(n125) );
	inv_0 U98 ( .x(n249), .a(A[3]) );
	inv_2 U99 ( .x(n338), .a(n61) );

endmodule


module EX_DW01_add_32_4_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n159, n160,
	n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
	n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
	n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
	n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
	n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
	n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
	n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
	n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
	n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
	n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
	n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
	n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
	n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
	n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
	n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
	n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
	n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n49,
	n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
	n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
	n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
	n92, n93, n94, n95, n96, n97, n98, n99;


	nand2i_2 U100 ( .x(n336), .a(n110), .b(n150) );
	nand2i_2 U101 ( .x(n285), .a(n110), .b(n148) );
	nand2i_2 U102 ( .x(n182), .a(n328), .b(n329) );
	inv_2 U103 ( .x(n222), .a(A[24]) );
	oai31_2 U104 ( .x(n261), .a(n98), .b(n110), .c(n100), .d(n262) );
	inv_2 U105 ( .x(n342), .a(n261) );
	inv_0 U106 ( .x(n224), .a(B[23]) );
	or3i_2 U107 ( .x(n255), .a(n148), .b(n224), .c(n110) );
	inv_2 U108 ( .x(n225), .a(A[23]) );
	or3i_2 U109 ( .x(n256), .a(n148), .b(n225), .c(n110) );
	inv_2 U11 ( .x(n58), .a(n60) );
	aoai211_1 U110 ( .x(n181), .a(n256), .b(n255), .c(n361), .d(n342) );
	inv_2 U111 ( .x(n281), .a(n329) );
	aoi21_1 U112 ( .x(n279), .a(n261), .b(n280), .c(n281) );
	inv_2 U113 ( .x(n344), .a(n255) );
	nand2i_2 U114 ( .x(n349), .a(n328), .b(n344) );
	inv_2 U115 ( .x(n343), .a(n256) );
	inv_2 U116 ( .x(n328), .a(n280) );
	nand2i_2 U117 ( .x(n350), .a(n328), .b(n343) );
	exor2_1 U118 ( .x(n180), .a(B[25]), .b(A[25]) );
	nor3i_2 U119 ( .x(n104), .a(n105), .b(n83), .c(n103) );
	nand2i_2 U12 ( .x(n264), .a(n127), .b(n232) );
	nand2_2 U120 ( .x(n105), .a(A[25]), .b(B[25]) );
	nor2i_3 U121 ( .x(n83), .a(B[25]), .b(n84) );
	exnor2_1 U122 ( .x(SUM[3]), .a(n174), .b(n106) );
	nor2i_1 U123 ( .x(n106), .a(n107), .b(n108) );
	exor2_1 U124 ( .x(SUM[2]), .a(n111), .b(n113) );
	exor2_1 U125 ( .x(SUM[6]), .a(n168), .b(n91) );
	nor2i_1 U126 ( .x(n91), .a(n50), .b(n67) );
	inv_2 U127 ( .x(n311), .a(n168) );
	exor2_1 U128 ( .x(SUM[12]), .a(n196), .b(n129) );
	oai21_1 U129 ( .x(n167), .a(n67), .b(n311), .c(n50) );
	inv_2 U13 ( .x(n254), .a(A[14]) );
	nor2i_1 U130 ( .x(n88), .a(n89), .b(n90) );
	inv_5 U131 ( .x(n90), .a(n273) );
	exor2_1 U132 ( .x(n178), .a(B[27]), .b(A[27]) );
	exor2_1 U133 ( .x(SUM[27]), .a(n71), .b(n178) );
	exor2_1 U134 ( .x(SUM[11]), .a(n197), .b(n132) );
	oai21_1 U135 ( .x(n197), .a(n137), .b(n338), .c(n136) );
	nor2i_1 U136 ( .x(n132), .a(n133), .b(n134) );
	inv_2 U137 ( .x(n134), .a(n242) );
	exor2_1 U138 ( .x(n187), .a(A[20]), .b(B[20]) );
	exor2_1 U139 ( .x(SUM[14]), .a(n194), .b(n123) );
	nor2_1 U14 ( .x(n102), .a(A[19]), .b(B[19]) );
	nand2i_2 U140 ( .x(n194), .a(n316), .b(n317) );
	nor2i_1 U141 ( .x(n123), .a(n124), .b(n125) );
	inv_2 U142 ( .x(n125), .a(n232) );
	inv_2 U143 ( .x(n318), .a(n194) );
	inv_2 U144 ( .x(n128), .a(n233) );
	nor2i_1 U145 ( .x(n126), .a(n127), .b(n128) );
	exor2_1 U146 ( .x(SUM[13]), .a(n195), .b(n126) );
	exor2_1 U147 ( .x(SUM[10]), .a(n198), .b(n135) );
	oai21_1 U148 ( .x(n198), .a(n164), .b(n87), .c(n86) );
	nor2i_0 U149 ( .x(n135), .a(n136), .b(n137) );
	oai211_1 U15 ( .x(n144), .a(n146), .b(n112), .c(n114), .d(n351) );
	inv_2 U150 ( .x(n338), .a(n198) );
	inv_2 U151 ( .x(n150), .a(n99) );
	aoi21_1 U152 ( .x(n147), .a(n148), .b(n149), .c(n150) );
	exnor2_1 U153 ( .x(n270), .a(A[22]), .b(B[22]) );
	aoi21_1 U154 ( .x(n109), .a(A[22]), .b(B[22]), .c(n110) );
	mux2i_1 U155 ( .x(SUM[22]), .d0(n109), .sl(n147), .d1(n270) );
	inv_2 U156 ( .x(n95), .a(n302) );
	nor2i_1 U157 ( .x(n93), .a(n94), .b(n95) );
	aoai211_1 U158 ( .x(n310), .a(n208), .b(n207), .c(n309), .d(n163) );
	exnor2_1 U159 ( .x(SUM[5]), .a(n169), .b(n93) );
	inv_0 U16 ( .x(n245), .a(A[10]) );
	exnor2_1 U160 ( .x(SUM[19]), .a(n116), .b(n188) );
	exor2_1 U161 ( .x(SUM[4]), .a(n170), .b(n162) );
	oai21_1 U162 ( .x(n170), .a(n108), .b(n174), .c(n107) );
	inv_2 U163 ( .x(n108), .a(n203) );
	inv_2 U164 ( .x(n174), .a(n293) );
	nor2i_1 U165 ( .x(n162), .a(n163), .b(n161) );
	inv_2 U166 ( .x(n309), .a(n170) );
	nand2i_2 U167 ( .x(n82), .a(n267), .b(n265) );
	exor2_1 U168 ( .x(n173), .a(B[30]), .b(A[30]) );
	exor2_1 U169 ( .x(n176), .a(A[28]), .b(B[28]) );
	nand2_2 U17 ( .x(n54), .a(n70), .b(n245) );
	inv_2 U170 ( .x(n219), .a(A[27]) );
	exnor2_1 U171 ( .x(SUM[28]), .a(n175), .b(n176) );
	exnor2_1 U172 ( .x(SUM[8]), .a(n165), .b(n166) );
	inv_2 U173 ( .x(n260), .a(A[30]) );
	exnor2_1 U175 ( .x(SUM[1]), .a(n357), .b(n354) );
	exnor2_1 U176 ( .x(SUM[9]), .a(n164), .b(n85) );
	inv_2 U177 ( .x(n164), .a(n308) );
	oai22_1 U178 ( .x(n308), .a(n214), .b(n215), .c(n240), .d(n307) );
	inv_2 U179 ( .x(n240), .a(n295) );
	inv_1 U18 ( .x(n70), .a(B[10]) );
	inv_2 U180 ( .x(n307), .a(n165) );
	nor2i_1 U181 ( .x(n85), .a(n86), .b(n87) );
	inv_2 U182 ( .x(n87), .a(n241) );
	exor2_1 U183 ( .x(SUM[15]), .a(n192), .b(n193) );
	exnor2_1 U184 ( .x(SUM[16]), .a(n191), .b(n120) );
	exor2_1 U186 ( .x(SUM[17]), .a(n189), .b(n190) );
	inv_2 U187 ( .x(n327), .a(n148) );
	nand2i_2 U188 ( .x(n185), .a(n327), .b(n99) );
	exnor2_1 U189 ( .x(SUM[21]), .a(n149), .b(n185) );
	nand3_3 U19 ( .x(n141), .a(n202), .b(n203), .c(n204) );
	exor2_1 U190 ( .x(SUM[23]), .a(n183), .b(n184) );
	exnor2_1 U191 ( .x(SUM[24]), .a(n181), .b(n182) );
	exnor2_1 U192 ( .x(SUM[25]), .a(n84), .b(n180) );
	inv_2 U193 ( .x(n74), .a(n73) );
	nand2_0 U194 ( .x(n50), .a(A[6]), .b(B[6]) );
	exnor2_1 U195 ( .x(n51), .a(B[29]), .b(A[29]) );
	or2_2 U196 ( .x(n52), .a(n145), .b(n105) );
	oa22_4 U197 ( .x(n53), .a(n57), .b(n252), .c(n124), .d(n58) );
	inv_2 U198 ( .x(n244), .a(n239) );
	oai21_1 U199 ( .x(n189), .a(n191), .b(n122), .c(n121) );
	or2_2 U20 ( .x(n62), .a(n160), .b(n107) );
	nand2i_4 U200 ( .x(n228), .a(n122), .b(n229) );
	inv_5 U201 ( .x(n122), .a(n320) );
	nand2i_0 U202 ( .x(n345), .a(A[5]), .b(n206) );
	nand2i_2 U203 ( .x(n233), .a(A[13]), .b(n253) );
	exnor2_1 U204 ( .x(SUM[20]), .a(n186), .b(n187) );
	oai211_1 U205 ( .x(n183), .a(n361), .b(n285), .c(n337), .d(n336) );
	oaoi211_1 U206 ( .x(n75), .a(B[20]), .b(A[20]), .c(n322), .d(n77) );
	nand2i_2 U207 ( .x(n302), .a(A[5]), .b(n206) );
	nand4_4 U208 ( .x(n210), .a(n59), .b(n211), .c(n212), .d(n213) );
	nor3i_5 U209 ( .x(n55), .a(n56), .b(n92), .c(n90) );
	nand2i_2 U21 ( .x(n319), .a(n65), .b(n195) );
	and2_1 U210 ( .x(n56), .a(B[5]), .b(A[5]) );
	nand2i_3 U211 ( .x(n273), .a(B[7]), .b(n205) );
	or2_8 U212 ( .x(n294), .a(A[6]), .b(B[6]) );
	inv_7 U213 ( .x(n92), .a(n294) );
	inv_1 U214 ( .x(n248), .a(A[17]) );
	nand2_0 U215 ( .x(n358), .a(n74), .b(A[1]) );
	nor2_1 U216 ( .x(n138), .a(n74), .b(A[1]) );
	nand2_2 U217 ( .x(n348), .a(n74), .b(A[1]) );
	nor2_1 U218 ( .x(n142), .a(n74), .b(A[1]) );
	nand2_1 U219 ( .x(n351), .a(B[1]), .b(A[1]) );
	nor2i_0 U22 ( .x(n96), .a(A[22]), .b(n97) );
	aoai211_4 U222 ( .x(n153), .a(n257), .b(n258), .c(n69), .d(n335) );
	inv_6 U223 ( .x(n69), .a(n353) );
	nand3i_2 U224 ( .x(n288), .a(n275), .b(n341), .c(n312) );
	nand2i_2 U225 ( .x(n341), .a(n86), .b(n54) );
	nor2_1 U226 ( .x(n160), .a(A[4]), .b(B[4]) );
	nor2_0 U227 ( .x(n161), .a(A[4]), .b(B[4]) );
	nand2_0 U228 ( .x(n163), .a(B[4]), .b(A[4]) );
	inv_12 U229 ( .x(n207), .a(A[4]) );
	nor2i_1 U23 ( .x(n98), .a(n99), .b(n96) );
	or2_1 U230 ( .x(n63), .a(A[5]), .b(B[5]) );
	inv_2 U231 ( .x(n206), .a(B[5]) );
	exor2_1 U232 ( .x(n193), .a(A[15]), .b(B[15]) );
	inv_2 U233 ( .x(n252), .a(B[15]) );
	inv_2 U234 ( .x(n246), .a(A[11]) );
	nand2_0 U235 ( .x(n274), .a(A[8]), .b(B[8]) );
	inv_0 U236 ( .x(n215), .a(A[8]) );
	inv_7 U237 ( .x(n205), .a(A[7]) );
	nand2_0 U238 ( .x(n89), .a(A[7]), .b(B[7]) );
	inv_0 U239 ( .x(n57), .a(A[15]) );
	inv_0 U24 ( .x(n304), .a(n112) );
	nand4_1 U240 ( .x(n177), .a(n333), .b(n332), .c(n331), .d(n52) );
	aoi23_1 U242 ( .x(n212), .a(A[7]), .b(B[7]), .c(A[6]), .d(B[6]), .e(n273) );
	nand2i_4 U243 ( .x(n232), .a(B[14]), .b(n254) );
	or2_2 U244 ( .x(n60), .a(A[15]), .b(B[15]) );
	and4i_5 U245 ( .x(n61), .a(n62), .b(n63), .c(n294), .d(n273) );
	nand3i_3 U246 ( .x(n230), .a(n231), .b(n232), .c(n233) );
	inv_2 U247 ( .x(n64), .a(n68) );
	inv_2 U249 ( .x(n157), .a(n284) );
	inv_2 U25 ( .x(n199), .a(A[2]) );
	nand2i_5 U250 ( .x(n352), .a(A[15]), .b(n252) );
	nand2i_2 U251 ( .x(n165), .a(n210), .b(n291) );
	oai21_1 U252 ( .x(n315), .a(n139), .b(n210), .c(n346) );
	nand3i_0 U253 ( .x(n65), .a(n231), .b(n232), .c(n233) );
	inv_10 U254 ( .x(n231), .a(n352) );
	inv_0 U255 ( .x(n66), .a(n92) );
	inv_2 U256 ( .x(n67), .a(n66) );
	aoai211_3 U257 ( .x(n79), .a(n350), .b(n349), .c(n76), .d(n279) );
	nand2_5 U259 ( .x(n114), .a(B[2]), .b(A[2]) );
	or3i_2 U26 ( .x(n306), .a(n301), .b(n201), .c(n200) );
	oai21_5 U260 ( .x(n263), .a(n231), .b(n264), .c(n53) );
	nand2i_2 U261 ( .x(n333), .a(n282), .b(n79) );
	nand2i_2 U262 ( .x(n332), .a(n283), .b(n79) );
	nor3i_2 U263 ( .x(n139), .a(n140), .b(n115), .c(n141) );
	aoi21_2 U265 ( .x(n151), .a(n152), .b(n153), .c(n154) );
	nor2_1 U266 ( .x(n101), .a(A[17]), .b(B[17]) );
	nand2_1 U267 ( .x(n298), .a(B[17]), .b(A[17]) );
	inv_4 U268 ( .x(n334), .a(n177) );
	inv_0 U269 ( .x(n71), .a(n334) );
	inv_2 U27 ( .x(n201), .a(n74) );
	nand2_1 U270 ( .x(n329), .a(A[24]), .b(B[24]) );
	nand2i_2 U271 ( .x(n320), .a(A[16]), .b(n247) );
	nand2_0 U272 ( .x(n94), .a(B[5]), .b(A[5]) );
	exnor2_3 U273 ( .x(SUM[31]), .a(n171), .b(n72) );
	inv_2 U274 ( .x(n72), .a(n172) );
	exor2_1 U275 ( .x(n172), .a(B[31]), .b(A[31]) );
	nor2i_0 U276 ( .x(n113), .a(n114), .b(n115) );
	inv_1 U277 ( .x(n303), .a(n114) );
	oai211_1 U278 ( .x(n140), .a(n142), .b(n112), .c(n114), .d(n348) );
	nand3i_1 U279 ( .x(n312), .a(n274), .b(n241), .c(n54) );
	aoi21_1 U28 ( .x(n111), .a(n112), .b(n358), .c(n356) );
	inv_0 U280 ( .x(n137), .a(n54) );
	nand4i_1 U281 ( .x(n239), .a(n240), .b(n54), .c(n241), .d(n242) );
	nand2_0 U282 ( .x(n354), .a(A[0]), .b(B[0]) );
	nor2_0 U283 ( .x(n355), .a(B[0]), .b(A[0]) );
	aoai211_2 U284 ( .x(n278), .a(B[18]), .b(A[18]), .c(n290), .d(n267) );
	nand2i_2 U285 ( .x(n280), .a(B[24]), .b(n222) );
	exor2_1 U286 ( .x(n190), .a(B[17]), .b(A[17]) );
	inv_3 U287 ( .x(n214), .a(B[8]) );
	ao21_1 U288 ( .x(n166), .a(A[8]), .b(B[8]), .c(n240) );
	inv_3 U289 ( .x(n216), .a(B[9]) );
	nand2_2 U29 ( .x(n112), .a(B[0]), .b(A[0]) );
	inv_2 U291 ( .x(n77), .a(n339) );
	inv_2 U292 ( .x(n78), .a(n226) );
	nand2_0 U293 ( .x(n339), .a(A[20]), .b(B[20]) );
	inv_0 U294 ( .x(n226), .a(B[20]) );
	inv_0 U295 ( .x(n186), .a(n322) );
	aoai211_1 U296 ( .x(n80), .a(n350), .b(n349), .c(n75), .d(n279) );
	nand4_1 U297 ( .x(n211), .a(n273), .b(n294), .c(n345), .d(n272) );
	nand2_0 U299 ( .x(n335), .a(B[28]), .b(A[28]) );
	inv_0 U30 ( .x(n227), .a(B[12]) );
	inv_0 U300 ( .x(n258), .a(B[28]) );
	inv_0 U301 ( .x(n257), .a(A[28]) );
	aoai211_3 U302 ( .x(n353), .a(n219), .b(n220), .c(n334), .d(n340) );
	nand2_2 U303 ( .x(n99), .a(B[21]), .b(A[21]) );
	nand2_1 U304 ( .x(n299), .a(B[16]), .b(A[16]) );
	nand2_0 U305 ( .x(n121), .a(B[16]), .b(A[16]) );
	exor2_3 U306 ( .x(SUM[7]), .a(n167), .b(n88) );
	exnor2_5 U308 ( .x(SUM[26]), .a(n104), .b(n179) );
	nand2_5 U309 ( .x(n107), .a(A[3]), .b(B[3]) );
	nand2i_0 U31 ( .x(n296), .a(A[12]), .b(n227) );
	nand2i_4 U310 ( .x(n234), .a(n235), .b(n236) );
	inv_6 U311 ( .x(n259), .a(B[30]) );
	exnor2_3 U312 ( .x(n268), .a(n359), .b(n249) );
	nor2_5 U313 ( .x(n202), .a(n92), .b(n90) );
	nor2i_5 U314 ( .x(n272), .a(B[4]), .b(n207) );
	nand2_2 U315 ( .x(n275), .a(n133), .b(n136) );
	oai21_4 U316 ( .x(n277), .a(n250), .b(n251), .c(n278) );
	nand2_2 U317 ( .x(n154), .a(n284), .b(n260) );
	exor2_3 U318 ( .x(n179), .a(A[26]), .b(B[26]) );
	nor2i_1 U32 ( .x(n129), .a(n130), .b(n131) );
	nand2i_4 U320 ( .x(n301), .a(B[2]), .b(n199) );
	nand2i_4 U321 ( .x(n203), .a(B[3]), .b(n209) );
	nand3i_3 U322 ( .x(n305), .a(n138), .b(n301), .c(n304) );
	nand3i_3 U323 ( .x(n293), .a(n303), .b(n306), .c(n305) );
	inv_5 U324 ( .x(n169), .a(n310) );
	oai21_4 U325 ( .x(n168), .a(n95), .b(n169), .c(n94) );
	nand2i_4 U326 ( .x(n242), .a(B[11]), .b(n246) );
	nand2i_4 U327 ( .x(n229), .a(B[17]), .b(n248) );
	nand2i_4 U328 ( .x(n321), .a(B[19]), .b(n251) );
	nand2i_4 U329 ( .x(n156), .a(B[29]), .b(n217) );
	nand2i_2 U33 ( .x(n314), .a(n134), .b(n288) );
	nand2_2 U330 ( .x(n337), .a(A[22]), .b(B[22]) );
	inv_5 U331 ( .x(n346), .a(n243) );
	nand2i_4 U332 ( .x(n326), .a(n130), .b(n347) );
	nand3i_3 U333 ( .x(n324), .a(n276), .b(n288), .c(n347) );
	aoai211_4 U334 ( .x(n323), .a(n238), .b(n263), .c(n277), .d(n321) );
	mux2i_3 U335 ( .x(n81), .d0(n271), .sl(B[18]), .d1(n268) );
	nand2_4 U336 ( .x(SUM[18]), .a(n81), .b(n82) );
	inv_6 U337 ( .x(n84), .a(n80) );
	inv_7 U338 ( .x(n110), .a(n300) );
	nand2i_6 U339 ( .x(n148), .a(A[21]), .b(n223) );
	inv_0 U34 ( .x(n292), .a(n141) );
	nor2i_5 U340 ( .x(n103), .a(A[25]), .b(n84) );
	nand2i_6 U341 ( .x(n241), .a(A[9]), .b(n216) );
	inv_10 U342 ( .x(n220), .a(B[27]) );
	inv_10 U343 ( .x(n208), .a(B[4]) );
	nor2_8 U344 ( .x(n100), .a(A[23]), .b(B[23]) );
	nand2_4 U345 ( .x(n262), .a(A[23]), .b(B[23]) );
	aoi21_4 U346 ( .x(n204), .a(n208), .b(n207), .c(n95) );
	aoi21_3 U347 ( .x(n359), .a(n118), .b(n236), .c(n360) );
	inv_3 U348 ( .x(n265), .a(n359) );
	inv_0 U349 ( .x(n360), .a(n266) );
	aoai211_1 U35 ( .x(n196), .a(n313), .b(n291), .c(n364), .d(n314) );
	inv_0 U350 ( .x(n191), .a(n118) );
	ao21_2 U351 ( .x(n266), .a(n298), .b(n299), .c(n101) );
	inv_5 U352 ( .x(n236), .a(n228) );
	nand2i_2 U353 ( .x(n118), .a(n263), .b(n319) );
	buf_3 U354 ( .x(n361), .a(n75) );
	inv_1 U355 ( .x(n175), .a(n353) );
	exnor2_3 U356 ( .x(SUM[29]), .a(n153), .b(n51) );
	nand4_4 U357 ( .x(n322), .a(n325), .b(n324), .c(n323), .d(n326) );
	oai211_3 U358 ( .x(n325), .a(n143), .b(n210), .c(n347), .d(n346) );
	ao21_3 U359 ( .x(n363), .a(n159), .b(n153), .c(n157) );
	nand2i_2 U36 ( .x(n330), .a(B[26]), .b(n221) );
	exnor2_3 U360 ( .x(SUM[30]), .a(n363), .b(n362) );
	inv_2 U361 ( .x(n362), .a(n173) );
	oai22_2 U362 ( .x(n171), .a(n155), .b(n260), .c(n151), .d(n259) );
	inv_0 U363 ( .x(n364), .a(n244) );
	aoi21_3 U364 ( .x(n155), .a(n156), .b(n153), .c(n157) );
	oaoi211_2 U365 ( .x(n76), .a(n78), .b(A[20]), .c(n322), .d(n77) );
	inv_2 U366 ( .x(n149), .a(n361) );
	inv_2 U37 ( .x(n221), .a(A[26]) );
	nand2_2 U38 ( .x(n331), .a(A[26]), .b(B[26]) );
	nand2i_2 U39 ( .x(n283), .a(n145), .b(A[25]) );
	nand2i_2 U40 ( .x(n282), .a(n145), .b(B[25]) );
	inv_2 U41 ( .x(n145), .a(n330) );
	nor2i_1 U42 ( .x(SUM[0]), .a(n354), .b(n355) );
	nand2_0 U43 ( .x(n133), .a(A[11]), .b(B[11]) );
	inv_5 U44 ( .x(n238), .a(n234) );
	inv_2 U45 ( .x(n251), .a(A[19]) );
	inv_0 U46 ( .x(n250), .a(B[19]) );
	nand2i_2 U47 ( .x(n276), .a(n131), .b(n242) );
	or3i_3 U48 ( .x(n237), .a(n238), .b(n102), .c(n230) );
	inv_5 U49 ( .x(n347), .a(n237) );
	nand2_2 U5 ( .x(n49), .a(n73), .b(n200) );
	nor3i_3 U50 ( .x(n143), .a(n144), .b(n115), .c(n141) );
	nand2_2 U51 ( .x(n195), .a(n287), .b(n315) );
	nand2_2 U52 ( .x(n317), .a(n195), .b(n233) );
	inv_0 U53 ( .x(n253), .a(B[13]) );
	inv_0 U54 ( .x(n316), .a(n127) );
	nand2_0 U55 ( .x(n127), .a(B[13]), .b(A[13]) );
	nand2i_2 U56 ( .x(n243), .a(n131), .b(n244) );
	inv_2 U57 ( .x(n115), .a(n301) );
	nand2_0 U58 ( .x(n130), .a(A[12]), .b(B[12]) );
	inv_2 U59 ( .x(n289), .a(n130) );
	inv_2 U6 ( .x(n146), .a(n49) );
	inv_2 U60 ( .x(n131), .a(n296) );
	nor2_1 U61 ( .x(n286), .a(n131), .b(n134) );
	aoi21_1 U62 ( .x(n287), .a(n286), .b(n288), .c(n289) );
	or2_2 U63 ( .x(n136), .a(n245), .b(n70) );
	inv_4 U64 ( .x(n97), .a(B[22]) );
	nand2i_2 U65 ( .x(n300), .a(A[22]), .b(n97) );
	exor2_1 U66 ( .x(n188), .a(A[19]), .b(B[19]) );
	inv_2 U67 ( .x(n290), .a(n266) );
	inv_0 U68 ( .x(n119), .a(n278) );
	nor2i_0 U69 ( .x(n117), .a(n267), .b(n228) );
	inv_10 U7 ( .x(n200), .a(A[1]) );
	aoi21_1 U70 ( .x(n116), .a(n117), .b(n118), .c(n119) );
	inv_0 U71 ( .x(n209), .a(A[3]) );
	nand2i_2 U72 ( .x(n267), .a(B[18]), .b(n249) );
	inv_7 U73 ( .x(n249), .a(A[18]) );
	inv_2 U74 ( .x(n235), .a(n267) );
	nor2i_1 U75 ( .x(n271), .a(A[18]), .b(n265) );
	nand2i_2 U77 ( .x(n159), .a(A[29]), .b(n218) );
	inv_2 U78 ( .x(n218), .a(B[29]) );
	nand2_2 U79 ( .x(n340), .a(B[27]), .b(A[27]) );
	inv_5 U8 ( .x(n73), .a(B[1]) );
	nand2i_2 U80 ( .x(n295), .a(A[8]), .b(n214) );
	nand2i_2 U81 ( .x(n152), .a(B[29]), .b(n217) );
	nand2_0 U82 ( .x(n284), .a(B[29]), .b(A[29]) );
	inv_2 U83 ( .x(n217), .a(A[29]) );
	nand2i_0 U84 ( .x(n297), .a(n74), .b(n200) );
	inv_2 U85 ( .x(n356), .a(n297) );
	nor2i_1 U86 ( .x(n357), .a(n358), .b(n356) );
	nand2_0 U87 ( .x(n86), .a(B[9]), .b(A[9]) );
	inv_0 U88 ( .x(n313), .a(n210) );
	nand2_2 U89 ( .x(n291), .a(n292), .b(n293) );
	inv_5 U90 ( .x(n213), .a(n55) );
	inv_4 U91 ( .x(n59), .a(n61) );
	inv_0 U92 ( .x(n68), .a(B[14]) );
	nand2i_2 U93 ( .x(n124), .a(n254), .b(n64) );
	oai21_1 U94 ( .x(n192), .a(n125), .b(n318), .c(n124) );
	nor2i_0 U95 ( .x(n120), .a(n121), .b(n122) );
	inv_3 U96 ( .x(n247), .a(B[16]) );
	inv_0 U98 ( .x(n223), .a(B[21]) );
	exor2_1 U99 ( .x(n184), .a(A[23]), .b(B[23]) );

endmodule


module EX_DW01_add_32_3_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n207, n208,
	n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
	n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
	n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
	n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
	n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
	n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
	n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
	n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
	n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
	n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
	n329, n330, n331, n332, n333, n335, n336, n337, n338, n339, n340, n341,
	n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
	n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
	n366, n367, n368, n369, n370, n371, n49, n50, n51, n52, n53, n54, n55,
	n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
	n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
	n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
	n98, n99;


	inv_2 U100 ( .x(n327), .a(n326) );
	oai21_1 U101 ( .x(n294), .a(A[2]), .b(B[2]), .c(n326) );
	aoi21_1 U102 ( .x(n144), .a(n145), .b(n369), .c(n146) );
	exnor2_1 U103 ( .x(SUM[2]), .a(n144), .b(n294) );
	oai21_1 U104 ( .x(n199), .a(n85), .b(n337), .c(n115) );
	exor2_1 U105 ( .x(SUM[6]), .a(n199), .b(n111) );
	exor2_1 U106 ( .x(SUM[12]), .a(n225), .b(n162) );
	nor2i_1 U107 ( .x(n162), .a(n163), .b(n164) );
	inv_2 U108 ( .x(n164), .a(n265) );
	inv_4 U109 ( .x(n340), .a(n225) );
	nor2_0 U11 ( .x(n77), .a(n127), .b(n78) );
	exor2_1 U110 ( .x(SUM[27]), .a(n91), .b(n209) );
	exor2_1 U111 ( .x(n209), .a(B[27]), .b(A[27]) );
	exnor2_1 U112 ( .x(SUM[11]), .a(n165), .b(n169) );
	exor2_1 U113 ( .x(n218), .a(A[20]), .b(B[20]) );
	inv_2 U114 ( .x(n354), .a(n223) );
	inv_4 U115 ( .x(n353), .a(n224) );
	inv_5 U116 ( .x(n161), .a(n55) );
	oai21_1 U117 ( .x(n223), .a(n161), .b(n353), .c(n160) );
	exor2_1 U118 ( .x(SUM[14]), .a(n223), .b(n156) );
	exor2_1 U119 ( .x(SUM[13]), .a(n224), .b(n159) );
	aoi21_2 U12 ( .x(n61), .a(n257), .b(n256), .c(n310) );
	exor2_1 U120 ( .x(SUM[10]), .a(n166), .b(n172) );
	inv_2 U121 ( .x(n190), .a(n122) );
	aoi21_1 U122 ( .x(n187), .a(n188), .b(n189), .c(n190) );
	exnor2_1 U123 ( .x(n297), .a(A[22]), .b(B[22]) );
	inv_5 U124 ( .x(n141), .a(n323) );
	aoi21_1 U125 ( .x(n140), .a(A[22]), .b(B[22]), .c(n141) );
	mux2i_1 U126 ( .x(SUM[22]), .d0(n140), .sl(n187), .d1(n297) );
	exor2_1 U127 ( .x(SUM[5]), .a(n200), .b(n114) );
	oai21_1 U128 ( .x(n200), .a(n118), .b(n336), .c(n64) );
	nor2i_0 U129 ( .x(n114), .a(n115), .b(n85) );
	nand2i_3 U13 ( .x(n267), .a(B[14]), .b(n261) );
	inv_0 U130 ( .x(n325), .a(n58) );
	inv_2 U131 ( .x(n337), .a(n200) );
	exor2_1 U132 ( .x(n219), .a(A[19]), .b(B[19]) );
	nor2i_1 U133 ( .x(n148), .a(n66), .b(n81) );
	oai21_1 U134 ( .x(n149), .a(n370), .b(n73), .c(n341) );
	aoi21_1 U135 ( .x(n71), .a(n289), .b(n285), .c(n125) );
	inv_0 U136 ( .x(n288), .a(n149) );
	exor2_1 U137 ( .x(SUM[4]), .a(n201), .b(n116) );
	inv_2 U138 ( .x(n139), .a(n324) );
	inv_2 U139 ( .x(n331), .a(n204) );
	inv_5 U14 ( .x(n158), .a(n267) );
	nor2i_1 U140 ( .x(n116), .a(n64), .b(n118) );
	inv_2 U141 ( .x(n118), .a(n234) );
	inv_2 U142 ( .x(n336), .a(n201) );
	nand2i_2 U143 ( .x(n105), .a(n66), .b(n287) );
	inv_0 U144 ( .x(n66), .a(n310) );
	inv_7 U145 ( .x(n126), .a(A[18]) );
	oai21_1 U146 ( .x(n287), .a(n288), .b(n81), .c(n49) );
	mux2i_1 U147 ( .x(n104), .d0(n298), .sl(B[18]), .d1(n295) );
	nor2i_0 U148 ( .x(n298), .a(A[18]), .b(n287) );
	exnor2_1 U149 ( .x(n295), .a(n296), .b(n126) );
	nor2_2 U15 ( .x(n304), .a(n161), .b(n163) );
	inv_2 U150 ( .x(n296), .a(n287) );
	exor2_1 U151 ( .x(n203), .a(B[30]), .b(A[30]) );
	inv_2 U152 ( .x(n194), .a(n279) );
	aoi21_1 U153 ( .x(n191), .a(n192), .b(n193), .c(n194) );
	exnor2_1 U156 ( .x(SUM[8]), .a(n196), .b(n197) );
	exor2_1 U157 ( .x(n205), .a(B[29]), .b(A[29]) );
	inv_0 U158 ( .x(n135), .a(B[30]) );
	inv_2 U159 ( .x(n244), .a(A[29]) );
	inv_2 U16 ( .x(n261), .a(A[14]) );
	exnor2_1 U160 ( .x(SUM[1]), .a(n368), .b(n365) );
	exnor2_1 U161 ( .x(SUM[9]), .a(n195), .b(n106) );
	inv_2 U162 ( .x(n195), .a(n335) );
	nor2i_1 U163 ( .x(n106), .a(n107), .b(n108) );
	inv_0 U164 ( .x(n108), .a(n272) );
	exor2_1 U165 ( .x(SUM[16]), .a(n149), .b(n154) );
	exnor2_1 U166 ( .x(SUM[17]), .a(n151), .b(n220) );
	exnor2_1 U167 ( .x(SUM[21]), .a(n142), .b(n95) );
	exor2_1 U168 ( .x(SUM[23]), .a(n215), .b(n216) );
	exor2_1 U169 ( .x(n212), .a(B[25]), .b(A[25]) );
	nand2_2 U17 ( .x(n266), .a(n69), .b(n260) );
	exor2_1 U170 ( .x(n211), .a(A[26]), .b(B[26]) );
	inv_2 U171 ( .x(n346), .a(n186) );
	exnor2_1 U172 ( .x(SUM[19]), .a(n147), .b(n219) );
	nand2_2 U173 ( .x(SUM[18]), .a(n104), .b(n105) );
	oa21_1 U174 ( .x(n49), .a(n124), .b(n155), .c(n286) );
	nand2i_4 U175 ( .x(n289), .a(B[18]), .b(n126) );
	inv_4 U176 ( .x(n310), .a(n289) );
	exor2_1 U177 ( .x(n207), .a(A[28]), .b(B[28]) );
	inv_1 U178 ( .x(n74), .a(B[17]) );
	and4i_4 U179 ( .x(n80), .a(n174), .b(n320), .c(n271), .d(n272) );
	inv_4 U18 ( .x(n69), .a(A[13]) );
	oai211_2 U180 ( .x(n56), .a(n58), .b(n299), .c(n301), .d(n332) );
	or3i_4 U181 ( .x(n268), .a(n61), .b(n127), .c(n78) );
	nor2_3 U182 ( .x(n127), .a(A[17]), .b(B[17]) );
	nand4_1 U183 ( .x(n292), .a(n272), .b(n271), .c(n305), .d(n167) );
	nand2i_3 U184 ( .x(n272), .a(A[9]), .b(n243) );
	nand2_2 U185 ( .x(n117), .a(B[4]), .b(A[4]) );
	inv_0 U186 ( .x(n54), .a(n53) );
	nand2_0 U187 ( .x(n50), .a(n61), .b(n77) );
	aoai211_1 U188 ( .x(n311), .a(n54), .b(n256), .c(n71), .d(n312) );
	inv_0 U189 ( .x(n51), .a(n52) );
	inv_7 U190 ( .x(n59), .a(A[5]) );
	aoai211_4 U191 ( .x(n60), .a(n363), .b(n362), .c(n62), .d(n314) );
	nand2_5 U192 ( .x(n338), .a(n52), .b(n258) );
	inv_2 U193 ( .x(n255), .a(A[16]) );
	aoi31_3 U194 ( .x(n293), .a(n167), .b(n271), .c(n306), .d(n175) );
	and2_5 U195 ( .x(n175), .a(n271), .b(n70) );
	oai21_2 U196 ( .x(n221), .a(n158), .b(n354), .c(n157) );
	nor2i_1 U197 ( .x(n156), .a(n157), .b(n158) );
	inv_4 U198 ( .x(n228), .a(B[5]) );
	inv_0 U199 ( .x(n53), .a(n257) );
	nand2_2 U20 ( .x(n303), .a(A[0]), .b(B[0]) );
	nand2_1 U200 ( .x(n112), .a(A[6]), .b(B[6]) );
	nand4i_2 U201 ( .x(n232), .a(n58), .b(n300), .c(n234), .d(n233) );
	and2_3 U202 ( .x(n301), .a(n112), .b(n57) );
	inv_2 U203 ( .x(n57), .a(n302) );
	or3i_4 U204 ( .x(n309), .a(n322), .b(n177), .c(n158) );
	aoai211_5 U206 ( .x(n84), .a(n246), .b(n247), .c(n349), .d(n356) );
	oaoi211_4 U207 ( .x(n62), .a(n98), .b(n97), .c(n217), .d(n96) );
	exor2_1 U208 ( .x(n222), .a(n51), .b(B[15]) );
	nand2_0 U209 ( .x(n308), .a(A[15]), .b(B[15]) );
	aoi22_1 U21 ( .x(n233), .a(n88), .b(n227), .c(n68), .d(n230) );
	inv_2 U210 ( .x(n258), .a(B[15]) );
	nand4i_3 U212 ( .x(n217), .a(n311), .b(n313), .c(n343), .d(n342) );
	nor2_4 U213 ( .x(n313), .a(n179), .b(n182) );
	and4i_4 U214 ( .x(n179), .a(n181), .b(n237), .c(n329), .d(n86) );
	inv_2 U215 ( .x(n68), .a(B[3]) );
	inv_0 U216 ( .x(n63), .a(n117) );
	inv_2 U217 ( .x(n64), .a(n63) );
	nand3i_0 U218 ( .x(n290), .a(n291), .b(n292), .c(n293) );
	inv_2 U219 ( .x(n339), .a(n290) );
	inv_4 U22 ( .x(n88), .a(B[7]) );
	nand2i_0 U220 ( .x(n324), .a(B[3]), .b(n230) );
	nor2i_2 U221 ( .x(n305), .a(A[8]), .b(n241) );
	inv_0 U222 ( .x(n242), .a(A[8]) );
	nand2i_6 U223 ( .x(n181), .a(n273), .b(n274) );
	inv_0 U224 ( .x(n67), .a(n75) );
	aoai211_2 U225 ( .x(n285), .a(n74), .b(n75), .c(n155), .d(n286) );
	inv_2 U226 ( .x(n256), .a(B[19]) );
	inv_2 U227 ( .x(n70), .a(n173) );
	nand2i_5 U228 ( .x(n300), .a(B[6]), .b(n226) );
	exor2_1 U229 ( .x(n220), .a(n67), .b(B[17]) );
	nor2i_1 U23 ( .x(n121), .a(n122), .b(n119) );
	nor2_0 U230 ( .x(n124), .a(B[17]), .b(n67) );
	or3i_4 U231 ( .x(n307), .a(n304), .b(n158), .c(n177) );
	nor2i_0 U232 ( .x(n137), .a(n138), .b(n139) );
	oai21_1 U233 ( .x(n201), .a(n139), .b(n331), .c(n138) );
	nand3_2 U234 ( .x(n283), .a(n307), .b(n309), .c(n308) );
	nor2_3 U235 ( .x(n182), .a(n181), .b(n183) );
	inv_0 U236 ( .x(n150), .a(n71) );
	nor2i_0 U237 ( .x(n172), .a(n173), .b(n174) );
	aoi21_1 U238 ( .x(n147), .a(n148), .b(n149), .c(n150) );
	nor2_1 U239 ( .x(n184), .a(n185), .b(n186) );
	nand2i_0 U24 ( .x(n330), .a(A[2]), .b(n238) );
	oai22_1 U240 ( .x(n335), .a(n241), .b(n242), .c(n270), .d(n370) );
	oai21_3 U241 ( .x(n225), .a(n370), .b(n269), .c(n339) );
	inv_0 U242 ( .x(n72), .a(n273) );
	inv_2 U243 ( .x(n73), .a(n72) );
	or3i_4 U244 ( .x(n282), .a(n284), .b(n176), .c(n283) );
	nand2i_2 U245 ( .x(n284), .a(n264), .b(n65) );
	or3i_2 U247 ( .x(n348), .a(n60), .b(n185), .c(n76) );
	inv_0 U248 ( .x(n76), .a(B[25]) );
	inv_0 U249 ( .x(n341), .a(n282) );
	inv_0 U25 ( .x(n238), .a(B[2]) );
	and2_3 U250 ( .x(n78), .a(n79), .b(n255) );
	inv_2 U251 ( .x(n79), .a(B[16]) );
	inv_4 U252 ( .x(n236), .a(n329) );
	ao21_1 U253 ( .x(n204), .a(n329), .b(n330), .c(n327) );
	oai21_5 U254 ( .x(n329), .a(n146), .b(n303), .c(n369) );
	nand2i_2 U255 ( .x(n363), .a(n344), .b(n358) );
	nand3i_1 U256 ( .x(n210), .a(n346), .b(n319), .c(n345) );
	nand2_4 U258 ( .x(n107), .a(B[9]), .b(A[9]) );
	inv_0 U259 ( .x(n269), .a(n80) );
	nand2_0 U26 ( .x(n326), .a(A[2]), .b(B[2]) );
	inv_0 U260 ( .x(n270), .a(n320) );
	nand2i_4 U261 ( .x(n167), .a(A[10]), .b(n263) );
	nand2i_8 U262 ( .x(n271), .a(A[11]), .b(n262) );
	nor2i_1 U263 ( .x(n154), .a(n155), .b(n78) );
	inv_2 U264 ( .x(n153), .a(n155) );
	inv_2 U265 ( .x(n185), .a(n347) );
	ao21_6 U266 ( .x(n90), .a(A[30]), .b(n99), .c(n132) );
	inv_1 U267 ( .x(n93), .a(n92) );
	aoi21_3 U268 ( .x(n132), .a(n133), .b(n134), .c(n135) );
	inv_7 U269 ( .x(n349), .a(n208) );
	inv_2 U27 ( .x(n231), .a(B[1]) );
	nand2i_0 U270 ( .x(n81), .a(n127), .b(n152) );
	inv_0 U271 ( .x(n82), .a(n217) );
	inv_2 U272 ( .x(n83), .a(n82) );
	inv_0 U274 ( .x(n85), .a(n325) );
	aoi21_2 U275 ( .x(n317), .a(n60), .b(n316), .c(n184) );
	nand3i_3 U276 ( .x(n208), .a(n130), .b(n348), .c(n317) );
	nand2i_4 U277 ( .x(n183), .a(n87), .b(n56) );
	nand2i_2 U278 ( .x(n315), .a(B[24]), .b(n249) );
	exor2_1 U279 ( .x(n214), .a(A[24]), .b(B[24]) );
	nand2_0 U28 ( .x(n145), .a(B[0]), .b(A[0]) );
	exor2_1 U280 ( .x(SUM[20]), .a(n83), .b(n218) );
	nand2i_4 U281 ( .x(n239), .a(n238), .b(n237) );
	nand2i_4 U282 ( .x(n235), .a(n236), .b(n237) );
	inv_5 U283 ( .x(n241), .a(B[8]) );
	ao21_1 U284 ( .x(n197), .a(A[8]), .b(B[8]), .c(n270) );
	inv_2 U286 ( .x(n86), .a(n180) );
	nor2_0 U287 ( .x(n180), .a(A[2]), .b(B[2]) );
	inv_3 U288 ( .x(n243), .a(B[9]) );
	nor2i_0 U289 ( .x(n109), .a(n110), .b(n87) );
	nand2_0 U29 ( .x(n170), .a(A[11]), .b(B[11]) );
	exnor2_5 U290 ( .x(SUM[31]), .a(n90), .b(n89) );
	inv_2 U291 ( .x(n89), .a(n202) );
	exor2_1 U292 ( .x(n202), .a(B[31]), .b(A[31]) );
	nand3i_0 U293 ( .x(n91), .a(n130), .b(n348), .c(n317) );
	inv_0 U294 ( .x(n92), .a(n60) );
	inv_0 U295 ( .x(n94), .a(n62) );
	inv_2 U296 ( .x(n95), .a(n94) );
	inv_0 U297 ( .x(n189), .a(n95) );
	inv_2 U298 ( .x(n98), .a(n253) );
	nand2_0 U299 ( .x(n355), .a(A[20]), .b(B[20]) );
	nand2_2 U30 ( .x(n110), .a(A[7]), .b(B[7]) );
	inv_0 U300 ( .x(n254), .a(A[20]) );
	inv_0 U301 ( .x(n253), .a(B[20]) );
	nand2_2 U302 ( .x(n122), .a(B[21]), .b(A[21]) );
	aoai211_1 U303 ( .x(n99), .a(n244), .b(n245), .c(n100), .d(n279) );
	nand2_1 U304 ( .x(n155), .a(A[16]), .b(B[16]) );
	nand2_0 U306 ( .x(n157), .a(A[14]), .b(B[14]) );
	and3i_1 U307 ( .x(n176), .a(n177), .b(B[14]), .c(A[14]) );
	inv_2 U308 ( .x(n193), .a(n100) );
	inv_2 U309 ( .x(n101), .a(n350) );
	inv_3 U31 ( .x(n227), .a(A[7]) );
	inv_2 U310 ( .x(n102), .a(n278) );
	inv_2 U311 ( .x(n103), .a(n277) );
	nand2_0 U312 ( .x(n350), .a(B[28]), .b(A[28]) );
	inv_0 U313 ( .x(n278), .a(B[28]) );
	inv_0 U314 ( .x(n277), .a(A[28]) );
	nand2_2 U316 ( .x(n163), .a(A[12]), .b(B[12]) );
	exor2_1 U317 ( .x(SUM[25]), .a(n93), .b(n212) );
	nand2_0 U318 ( .x(n319), .a(B[25]), .b(n93) );
	nand2_0 U319 ( .x(n345), .a(A[25]), .b(n93) );
	nand2i_2 U32 ( .x(n347), .a(B[26]), .b(n248) );
	nor2i_0 U320 ( .x(n111), .a(n112), .b(n113) );
	inv_0 U321 ( .x(n321), .a(n112) );
	nand2_1 U322 ( .x(n173), .a(B[10]), .b(A[10]) );
	inv_6 U323 ( .x(n263), .a(B[10]) );
	exor2_3 U324 ( .x(SUM[7]), .a(n198), .b(n109) );
	exnor2_3 U325 ( .x(SUM[30]), .a(n191), .b(n203) );
	exnor2_3 U326 ( .x(SUM[28]), .a(n371), .b(n207) );
	exor2_3 U327 ( .x(SUM[26]), .a(n210), .b(n211) );
	exor2_3 U328 ( .x(SUM[15]), .a(n221), .b(n222) );
	inv_6 U329 ( .x(n251), .a(B[23]) );
	inv_2 U33 ( .x(n248), .a(A[26]) );
	inv_6 U330 ( .x(n134), .a(A[30]) );
	nand3i_3 U331 ( .x(n299), .a(n138), .b(n300), .c(n234) );
	nand2i_4 U332 ( .x(n328), .a(A[1]), .b(n231) );
	inv_5 U333 ( .x(n146), .a(n328) );
	ao211_5 U334 ( .x(n332), .a(n117), .b(n115), .c(n58), .d(n113) );
	ao21_4 U335 ( .x(n198), .a(n199), .b(n300), .c(n321) );
	nand2_2 U336 ( .x(n352), .a(A[22]), .b(B[22]) );
	oai21_4 U337 ( .x(n224), .a(n340), .b(n164), .c(n163) );
	inv_5 U338 ( .x(n358), .a(n276) );
	nand2i_4 U339 ( .x(n342), .a(n50), .b(n282) );
	nor2i_1 U34 ( .x(n130), .a(A[26]), .b(n131) );
	nand3i_5 U340 ( .x(n343), .a(n240), .b(n360), .c(n361) );
	nand2i_6 U341 ( .x(n188), .a(A[21]), .b(n250) );
	or3i_5 U342 ( .x(n276), .a(n188), .b(n252), .c(n141) );
	or3i_5 U343 ( .x(n275), .a(n188), .b(n251), .c(n141) );
	inv_6 U344 ( .x(n113), .a(n300) );
	nand2i_6 U345 ( .x(n323), .a(A[22]), .b(n120) );
	nor2i_5 U346 ( .x(n316), .a(A[25]), .b(n185) );
	inv_10 U347 ( .x(n246), .a(A[27]) );
	inv_10 U348 ( .x(n247), .a(B[27]) );
	nand2_4 U349 ( .x(n356), .a(B[27]), .b(A[27]) );
	inv_2 U35 ( .x(n131), .a(B[26]) );
	nand2i_6 U350 ( .x(n234), .a(A[4]), .b(n229) );
	inv_10 U351 ( .x(n262), .a(B[11]) );
	inv_6 U352 ( .x(n177), .a(n338) );
	inv_14 U353 ( .x(n120), .a(B[22]) );
	nor2_8 U354 ( .x(n123), .a(A[23]), .b(B[23]) );
	nand2_4 U355 ( .x(n281), .a(A[23]), .b(B[23]) );
	inv_10 U356 ( .x(n229), .a(B[4]) );
	nor2i_8 U357 ( .x(n119), .a(A[22]), .b(n120) );
	oa222_4 U358 ( .x(n370), .a(n239), .b(n240), .c(n87), .d(n333), .e(n178),
		.f(n235) );
	inv_0 U359 ( .x(n196), .a(n370) );
	nor2i_1 U36 ( .x(SUM[0]), .a(n365), .b(n366) );
	inv_3 U360 ( .x(n333), .a(n56) );
	inv_0 U361 ( .x(n240), .a(A[2]) );
	aoi221_4 U362 ( .x(n100), .a(n103), .b(n364), .c(n84), .d(n102), .e(n101) );
	aoai211_4 U363 ( .x(n364), .a(n246), .b(n247), .c(n349), .d(n356) );
	inv_5 U364 ( .x(n133), .a(n136) );
	aoai211_4 U365 ( .x(n136), .a(n244), .b(n245), .c(n100), .d(n279) );
	inv_3 U366 ( .x(n361), .a(n181) );
	exnor2_2 U367 ( .x(SUM[29]), .a(n100), .b(n205) );
	inv_2 U368 ( .x(n371), .a(n364) );
	nand4_3 U369 ( .x(n264), .a(n338), .b(n265), .c(n266), .d(n267) );
	nor2_1 U37 ( .x(n366), .a(B[0]), .b(A[0]) );
	nand2i_4 U370 ( .x(n265), .a(B[12]), .b(n259) );
	nand2i_4 U371 ( .x(n273), .a(n264), .b(n80) );
	inv_4 U372 ( .x(n260), .a(B[13]) );
	inv_2 U38 ( .x(n291), .a(n170) );
	inv_2 U39 ( .x(n171), .a(n271) );
	nor2i_1 U40 ( .x(n169), .a(n170), .b(n171) );
	aoi21_1 U41 ( .x(n165), .a(n166), .b(n167), .c(n168) );
	inv_4 U42 ( .x(n274), .a(n268) );
	inv_5 U43 ( .x(n257), .a(A[19]) );
	nand2_0 U44 ( .x(n312), .a(A[19]), .b(B[19]) );
	nor2i_1 U45 ( .x(n159), .a(n160), .b(n161) );
	nand2_1 U46 ( .x(n160), .a(B[13]), .b(A[13]) );
	nand2_2 U47 ( .x(n55), .a(n69), .b(n260) );
	inv_2 U48 ( .x(n322), .a(n160) );
	inv_2 U49 ( .x(n259), .a(A[12]) );
	nand2i_4 U5 ( .x(n320), .a(A[8]), .b(n241) );
	inv_0 U50 ( .x(n168), .a(n173) );
	oai21_1 U51 ( .x(n166), .a(n195), .b(n108), .c(n107) );
	nand2_1 U52 ( .x(n115), .a(B[5]), .b(A[5]) );
	and2_1 U53 ( .x(n125), .a(B[18]), .b(A[18]) );
	inv_5 U54 ( .x(n75), .a(A[17]) );
	inv_2 U55 ( .x(n174), .a(n167) );
	inv_2 U56 ( .x(n230), .a(A[3]) );
	nand2_2 U57 ( .x(n138), .a(A[3]), .b(B[3]) );
	nand2_2 U58 ( .x(n286), .a(A[17]), .b(B[17]) );
	nand2i_2 U59 ( .x(n192), .a(A[29]), .b(n245) );
	inv_5 U6 ( .x(n226), .a(A[6]) );
	and2_6 U60 ( .x(n58), .a(n59), .b(n228) );
	inv_2 U61 ( .x(n302), .a(n110) );
	inv_5 U62 ( .x(n237), .a(n232) );
	nor2_0 U63 ( .x(n178), .a(A[2]), .b(B[2]) );
	and2_1 U64 ( .x(n87), .a(n88), .b(n227) );
	inv_5 U65 ( .x(n360), .a(n239) );
	inv_2 U66 ( .x(n245), .a(B[29]) );
	nand2_2 U68 ( .x(n279), .a(B[29]), .b(A[29]) );
	nand2_0 U69 ( .x(n365), .a(A[0]), .b(B[0]) );
	nand3i_2 U7 ( .x(n65), .a(n291), .b(n292), .c(n293) );
	nor2_1 U70 ( .x(n367), .a(B[1]), .b(A[1]) );
	nand2_2 U71 ( .x(n369), .a(B[1]), .b(A[1]) );
	nor2i_1 U72 ( .x(n368), .a(n369), .b(n367) );
	inv_2 U73 ( .x(n306), .a(n107) );
	inv_2 U75 ( .x(n152), .a(n78) );
	aoi21_1 U76 ( .x(n151), .a(n152), .b(n149), .c(n153) );
	inv_0 U77 ( .x(n250), .a(B[21]) );
	inv_2 U78 ( .x(n143), .a(n188) );
	nor2i_1 U79 ( .x(n142), .a(n122), .b(n143) );
	inv_10 U8 ( .x(n52), .a(A[15]) );
	exor2_1 U80 ( .x(n216), .a(A[23]), .b(B[23]) );
	nand2i_0 U81 ( .x(n351), .a(n141), .b(n190) );
	nand2i_2 U82 ( .x(n318), .a(n141), .b(n188) );
	oai211_1 U83 ( .x(n215), .a(n95), .b(n318), .c(n352), .d(n351) );
	exor2_1 U84 ( .x(SUM[24]), .a(n213), .b(n214) );
	aoai211_1 U85 ( .x(n213), .a(n276), .b(n275), .c(n95), .d(n357) );
	aoi21_1 U86 ( .x(n314), .a(n280), .b(n315), .c(n128) );
	oai31_1 U87 ( .x(n280), .a(n121), .b(n141), .c(n123), .d(n281) );
	nor2i_1 U88 ( .x(n128), .a(A[24]), .b(n129) );
	inv_2 U89 ( .x(n129), .a(B[24]) );
	inv_2 U90 ( .x(n357), .a(n280) );
	inv_2 U91 ( .x(n96), .a(n355) );
	inv_2 U92 ( .x(n97), .a(n254) );
	nand2i_2 U93 ( .x(n362), .a(n344), .b(n359) );
	inv_2 U94 ( .x(n359), .a(n275) );
	inv_2 U95 ( .x(n344), .a(n315) );
	inv_2 U96 ( .x(n249), .a(A[24]) );
	inv_2 U97 ( .x(n252), .a(A[23]) );
	nand2_2 U98 ( .x(n186), .a(A[25]), .b(B[25]) );
	exor2_1 U99 ( .x(SUM[3]), .a(n204), .b(n137) );

endmodule


module EX_DW01_add_32_7_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n190, n191, n192, n193, n194, n195, n197,
	n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
	n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
	n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
	n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
	n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
	n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
	n270, n271, n272, n273, n275, n276, n277, n278, n279, n280, n281, n282,
	n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
	n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
	n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
	n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
	n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
	n343, n344, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
	n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
	n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
	n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	inv_2 U10 ( .x(n60), .a(B[14]) );
	inv_2 U100 ( .x(n331), .a(n267) );
	or3i_2 U101 ( .x(n267), .a(n190), .b(n245), .c(n138) );
	inv_2 U102 ( .x(n245), .a(B[23]) );
	nand2i_2 U103 ( .x(n333), .a(n322), .b(n330) );
	inv_2 U104 ( .x(n322), .a(n295) );
	nand2i_0 U105 ( .x(n295), .a(B[24]), .b(n242) );
	inv_2 U106 ( .x(n242), .a(A[24]) );
	inv_2 U107 ( .x(n330), .a(n268) );
	or3i_2 U108 ( .x(n268), .a(n190), .b(n246), .c(n138) );
	inv_2 U109 ( .x(n246), .a(A[23]) );
	nor2_0 U11 ( .x(n336), .a(B[0]), .b(A[0]) );
	nand2_2 U110 ( .x(n184), .a(n55), .b(B[25]) );
	exor2_1 U111 ( .x(SUM[3]), .a(n203), .b(n134) );
	inv_2 U112 ( .x(n309), .a(n308) );
	nor2i_1 U113 ( .x(n134), .a(n135), .b(n136) );
	inv_2 U114 ( .x(n136), .a(n306) );
	inv_2 U115 ( .x(n313), .a(n203) );
	exnor2_1 U116 ( .x(SUM[2]), .a(n139), .b(n277) );
	exor2_1 U117 ( .x(SUM[6]), .a(n200), .b(n107) );
	exnor2_1 U118 ( .x(SUM[12]), .a(n50), .b(n157) );
	nor2i_0 U119 ( .x(n157), .a(n158), .b(n159) );
	nor2_1 U12 ( .x(n121), .a(A[17]), .b(B[17]) );
	inv_0 U120 ( .x(n159), .a(n251) );
	exor2_1 U121 ( .x(n207), .a(B[27]), .b(A[27]) );
	exnor2_1 U122 ( .x(SUM[11]), .a(n160), .b(n164) );
	inv_2 U123 ( .x(n163), .a(n168) );
	nor2i_1 U124 ( .x(n164), .a(n165), .b(n166) );
	exor2_1 U125 ( .x(n215), .a(n95), .b(B[20]) );
	exnor2_1 U126 ( .x(SUM[20]), .a(n89), .b(n215) );
	exor2_1 U127 ( .x(SUM[14]), .a(n220), .b(n151) );
	exor2_1 U128 ( .x(SUM[13]), .a(n221), .b(n154) );
	exor2_1 U129 ( .x(SUM[10]), .a(n161), .b(n167) );
	nand2i_2 U13 ( .x(n323), .a(B[26]), .b(n241) );
	oai21_1 U130 ( .x(n161), .a(n49), .b(n103), .c(n102) );
	nor2i_1 U131 ( .x(n167), .a(n168), .b(n169) );
	inv_0 U132 ( .x(n169), .a(n162) );
	inv_2 U133 ( .x(n191), .a(n118) );
	exnor2_1 U134 ( .x(n280), .a(A[22]), .b(B[22]) );
	aoi21_1 U135 ( .x(n137), .a(A[22]), .b(B[22]), .c(n138) );
	exor2_1 U137 ( .x(SUM[5]), .a(n201), .b(n109) );
	exnor2_1 U138 ( .x(SUM[19]), .a(n142), .b(n216) );
	exor2_1 U139 ( .x(n216), .a(A[19]), .b(B[19]) );
	inv_2 U14 ( .x(n241), .a(A[26]) );
	inv_2 U140 ( .x(n114), .a(n229) );
	nor2i_1 U141 ( .x(n112), .a(n113), .b(n114) );
	exor2_1 U142 ( .x(SUM[4]), .a(n202), .b(n112) );
	nand2i_0 U143 ( .x(n100), .a(n276), .b(n273) );
	exnor2_1 U144 ( .x(SUM[28]), .a(n204), .b(n205) );
	exnor2_1 U145 ( .x(SUM[8]), .a(n197), .b(n198) );
	inv_5 U146 ( .x(n235), .a(A[2]) );
	inv_5 U147 ( .x(n106), .a(n305) );
	inv_0 U149 ( .x(n132), .a(B[30]) );
	and2_3 U15 ( .x(n81), .a(A[0]), .b(B[0]) );
	inv_2 U150 ( .x(n131), .a(A[30]) );
	inv_5 U151 ( .x(n130), .a(n133) );
	inv_2 U152 ( .x(n239), .a(A[29]) );
	nor2i_1 U153 ( .x(n101), .a(n102), .b(n103) );
	exnor2_1 U154 ( .x(SUM[9]), .a(n49), .b(n101) );
	inv_5 U155 ( .x(n252), .a(n59) );
	oai21_1 U156 ( .x(n218), .a(n153), .b(n326), .c(n152) );
	exor2_2 U157 ( .x(SUM[15]), .a(n218), .b(n219) );
	exnor2_1 U158 ( .x(SUM[17]), .a(n145), .b(n217) );
	inv_2 U159 ( .x(n301), .a(n190) );
	nor2i_3 U16 ( .x(n69), .a(n98), .b(A[6]) );
	nand2i_2 U160 ( .x(n214), .a(n301), .b(n118) );
	inv_2 U161 ( .x(n94), .a(n327) );
	inv_1 U162 ( .x(n247), .a(B[20]) );
	exnor2_1 U163 ( .x(SUM[23]), .a(n185), .b(n213) );
	exor2_1 U164 ( .x(n213), .a(A[23]), .b(B[23]) );
	exnor2_1 U165 ( .x(SUM[25]), .a(n210), .b(n211) );
	exor2_1 U166 ( .x(n211), .a(B[25]), .b(n55) );
	exor2_1 U167 ( .x(n209), .a(A[26]), .b(B[26]) );
	inv_2 U168 ( .x(n269), .a(B[25]) );
	inv_5 U169 ( .x(n210), .a(n299) );
	nor2_2 U17 ( .x(n228), .a(n106), .b(n136) );
	oai221_1 U170 ( .x(n208), .a(n210), .b(n269), .c(n210), .d(n54), .e(n184) );
	exor2_1 U171 ( .x(SUM[26]), .a(n208), .b(n209) );
	ao21_2 U173 ( .x(n88), .a(n133), .b(A[30]), .c(n129) );
	inv_2 U174 ( .x(n293), .a(n82) );
	oa22_1 U175 ( .x(n49), .a(n236), .b(n237), .c(n253), .d(n316) );
	aoi22_1 U176 ( .x(n50), .a(n329), .b(n255), .c(n197), .d(n73) );
	inv_2 U177 ( .x(n55), .a(n54) );
	inv_2 U178 ( .x(n54), .a(A[25]) );
	inv_1 U179 ( .x(n86), .a(B[19]) );
	nand2i_2 U18 ( .x(n306), .a(B[3]), .b(n225) );
	exnor2_1 U180 ( .x(n51), .a(B[31]), .b(A[31]) );
	inv_2 U181 ( .x(n174), .a(n258) );
	nand2i_2 U182 ( .x(n258), .a(n75), .b(n259) );
	exnor2_1 U183 ( .x(n52), .a(B[30]), .b(A[30]) );
	exnor2_1 U184 ( .x(n53), .a(B[29]), .b(A[29]) );
	exor2_1 U186 ( .x(n205), .a(A[28]), .b(B[28]) );
	inv_2 U187 ( .x(n95), .a(n248) );
	oai211_2 U188 ( .x(n291), .a(n156), .b(n158), .c(n155), .d(n152) );
	nand2_2 U189 ( .x(n158), .a(A[12]), .b(B[12]) );
	inv_2 U19 ( .x(n225), .a(A[3]) );
	nand2i_2 U190 ( .x(n307), .a(A[5]), .b(n223) );
	nand2_1 U191 ( .x(n110), .a(B[5]), .b(A[5]) );
	nor2i_5 U192 ( .x(n97), .a(A[6]), .b(n98) );
	ao211_5 U193 ( .x(n314), .a(n113), .b(n110), .c(n111), .d(n69) );
	nor2_6 U194 ( .x(n176), .a(n177), .b(n178) );
	nor2i_0 U195 ( .x(n143), .a(n276), .b(n249) );
	oai21_1 U196 ( .x(n273), .a(n340), .b(n249), .c(n275) );
	nor2_0 U197 ( .x(n337), .a(n85), .b(A[1]) );
	nand2i_2 U198 ( .x(n310), .a(A[1]), .b(n226) );
	inv_2 U199 ( .x(n79), .a(A[1]) );
	nand2_2 U20 ( .x(n335), .a(A[0]), .b(B[0]) );
	nand2_3 U200 ( .x(n135), .a(A[3]), .b(B[3]) );
	nor2_2 U201 ( .x(n230), .a(n111), .b(n69) );
	oai21_2 U202 ( .x(n200), .a(n111), .b(n318), .c(n110) );
	inv_8 U203 ( .x(n111), .a(n307) );
	aoi21_1 U204 ( .x(n142), .a(n143), .b(n144), .c(n82) );
	aoi21_1 U205 ( .x(n145), .a(n146), .b(n144), .c(n147) );
	exor2_1 U206 ( .x(SUM[16]), .a(n144), .b(n148) );
	exnor2_1 U208 ( .x(SUM[21]), .a(n92), .b(n214) );
	nor2i_1 U21 ( .x(n338), .a(n339), .b(n337) );
	aoi21_1 U210 ( .x(n185), .a(n186), .b(n92), .c(n188) );
	aoi21_1 U211 ( .x(n192), .a(n193), .b(n92), .c(n194) );
	inv_0 U212 ( .x(n187), .a(n93) );
	ao23_3 U214 ( .x(n63), .a(B[15]), .b(A[15]), .c(n291), .d(n252), .e(n70) );
	nand4_1 U215 ( .x(n250), .a(n252), .b(n319), .c(n251), .d(n70) );
	nand2_2 U216 ( .x(n113), .a(B[4]), .b(A[4]) );
	nand2i_2 U217 ( .x(n229), .a(A[4]), .b(n224) );
	inv_2 U218 ( .x(n223), .a(B[5]) );
	inv_2 U219 ( .x(n56), .a(n170) );
	inv_2 U22 ( .x(n62), .a(n166) );
	oai222_4 U220 ( .x(n321), .a(n235), .b(n288), .c(n179), .d(n122), .e(n181),
		.f(n286) );
	exor2_1 U221 ( .x(n219), .a(A[15]), .b(B[15]) );
	inv_5 U222 ( .x(n71), .a(B[15]) );
	and4_5 U223 ( .x(n73), .a(n303), .b(n254), .c(n162), .d(n255) );
	nand2_2 U224 ( .x(n165), .a(A[11]), .b(B[11]) );
	nand2i_2 U225 ( .x(n303), .a(A[8]), .b(n236) );
	inv_0 U226 ( .x(n237), .a(A[8]) );
	ao21_1 U227 ( .x(n198), .a(A[8]), .b(B[8]), .c(n253) );
	nand2_1 U228 ( .x(n289), .a(A[8]), .b(B[8]) );
	nand2_1 U229 ( .x(n105), .a(A[7]), .b(B[7]) );
	inv_5 U23 ( .x(n173), .a(n74) );
	and4i_2 U231 ( .x(n58), .a(n59), .b(n319), .c(n251), .d(n70) );
	nand2i_2 U232 ( .x(n251), .a(B[12]), .b(n264) );
	inv_2 U233 ( .x(n65), .a(A[6]) );
	exnor2_3 U234 ( .x(SUM[30]), .a(n61), .b(n52) );
	oai21_1 U235 ( .x(n61), .a(n57), .b(n64), .c(n270) );
	ao31_6 U236 ( .x(n272), .a(n329), .b(n62), .c(n58), .d(n63) );
	inv_2 U237 ( .x(n64), .a(n195) );
	ao221_3 U238 ( .x(n282), .a(n98), .b(n65), .c(n66), .d(n224), .e(n135) );
	inv_5 U239 ( .x(n224), .a(B[4]) );
	nor2i_1 U24 ( .x(n123), .a(A[19]), .b(n86) );
	inv_10 U240 ( .x(n68), .a(A[13]) );
	inv_0 U241 ( .x(n253), .a(n303) );
	inv_2 U242 ( .x(n166), .a(n255) );
	exor2_1 U243 ( .x(SUM[27]), .a(n206), .b(n207) );
	nand2_5 U246 ( .x(n74), .a(n174), .b(n272) );
	inv_0 U247 ( .x(n175), .a(n272) );
	oai211_4 U248 ( .x(n292), .a(n282), .b(n111), .c(n284), .d(n314) );
	inv_0 U249 ( .x(n276), .a(n75) );
	nand2_2 U25 ( .x(n271), .a(A[23]), .b(B[23]) );
	inv_5 U250 ( .x(n76), .a(B[18]) );
	inv_16 U251 ( .x(n261), .a(A[18]) );
	inv_0 U253 ( .x(n339), .a(n78) );
	inv_6 U254 ( .x(n80), .a(B[1]) );
	inv_0 U255 ( .x(n141), .a(n310) );
	nand2_4 U256 ( .x(n102), .a(A[9]), .b(B[9]) );
	nor2_0 U257 ( .x(n120), .a(B[17]), .b(A[17]) );
	oaoi211_2 U258 ( .x(n82), .a(n83), .b(n261), .c(n275), .d(n75) );
	inv_0 U259 ( .x(n83), .a(B[18]) );
	nor2_1 U26 ( .x(n119), .a(A[23]), .b(B[23]) );
	ao21_3 U260 ( .x(n275), .a(n302), .b(n149), .c(n120) );
	inv_2 U261 ( .x(n260), .a(A[16]) );
	nand2_0 U262 ( .x(n302), .a(A[17]), .b(B[17]) );
	inv_2 U264 ( .x(n265), .a(A[10]) );
	inv_0 U265 ( .x(n84), .a(B[1]) );
	inv_2 U266 ( .x(n85), .a(n84) );
	ao211_5 U267 ( .x(n177), .a(n87), .b(n86), .c(n258), .d(n256) );
	inv_2 U268 ( .x(n87), .a(A[19]) );
	exnor2_3 U269 ( .x(SUM[31]), .a(n88), .b(n51) );
	nor2i_1 U27 ( .x(n117), .a(n118), .b(n115) );
	oa222_1 U270 ( .x(n89), .a(n235), .b(n288), .c(n179), .d(n122), .e(n181),
		.f(n286) );
	nand2i_5 U271 ( .x(n286), .a(n231), .b(n287) );
	nand2i_4 U272 ( .x(n288), .a(n234), .b(n287) );
	exor2_1 U273 ( .x(n212), .a(A[24]), .b(B[24]) );
	exor2_1 U274 ( .x(n217), .a(A[17]), .b(B[17]) );
	inv_2 U275 ( .x(n90), .a(n324) );
	inv_0 U276 ( .x(n204), .a(n334) );
	nand2_0 U277 ( .x(n324), .a(B[28]), .b(A[28]) );
	inv_2 U278 ( .x(n91), .a(n187) );
	inv_4 U279 ( .x(n92), .a(n91) );
	nor2i_1 U28 ( .x(n115), .a(A[22]), .b(n116) );
	inv_2 U280 ( .x(n96), .a(n247) );
	nand2_0 U281 ( .x(n327), .a(A[20]), .b(B[20]) );
	inv_0 U282 ( .x(n248), .a(A[20]) );
	nand2_3 U283 ( .x(n118), .a(B[21]), .b(A[21]) );
	aoi21_1 U284 ( .x(n160), .a(n161), .b(n162), .c(n163) );
	nand2i_3 U285 ( .x(n162), .a(B[10]), .b(n265) );
	nand2i_2 U286 ( .x(n305), .a(B[7]), .b(n222) );
	nand2_2 U287 ( .x(n168), .a(A[10]), .b(B[10]) );
	nor2i_5 U288 ( .x(n104), .a(n105), .b(n106) );
	nor2_5 U289 ( .x(n172), .a(A[2]), .b(B[2]) );
	inv_2 U29 ( .x(n116), .a(B[22]) );
	nor3_5 U290 ( .x(n179), .a(n176), .b(n173), .c(n180) );
	nor2_5 U291 ( .x(n181), .a(A[2]), .b(B[2]) );
	nor2_5 U292 ( .x(n182), .a(n183), .b(n184) );
	exor2_3 U293 ( .x(SUM[7]), .a(n199), .b(n104) );
	exnor2_3 U294 ( .x(SUM[24]), .a(n192), .b(n212) );
	inv_6 U295 ( .x(n240), .a(B[29]) );
	inv_6 U296 ( .x(n264), .a(A[12]) );
	exnor2_3 U297 ( .x(n278), .a(n279), .b(n261) );
	nor2i_5 U298 ( .x(n284), .a(n108), .b(n285) );
	nand2_2 U299 ( .x(n290), .a(n165), .b(n168) );
	nand2i_2 U30 ( .x(n312), .a(A[2]), .b(n233) );
	nand2i_4 U300 ( .x(n180), .a(n123), .b(n293) );
	aoi21_3 U301 ( .x(n298), .a(n296), .b(n299), .c(n126) );
	aoi21_3 U302 ( .x(n300), .a(n297), .b(n299), .c(n182) );
	nand2_5 U303 ( .x(n308), .a(A[2]), .b(B[2]) );
	ao21_4 U304 ( .x(n203), .a(n311), .b(n312), .c(n309) );
	oai222_4 U305 ( .x(n197), .a(n234), .b(n235), .c(n106), .d(n315), .e(n172),
		.f(n231) );
	oai21_4 U306 ( .x(n202), .a(n136), .b(n313), .c(n135) );
	inv_5 U307 ( .x(n317), .a(n202) );
	oai21_4 U308 ( .x(n201), .a(n114), .b(n317), .c(n113) );
	inv_5 U309 ( .x(n318), .a(n201) );
	oai21_1 U31 ( .x(n277), .a(A[2]), .b(B[2]), .c(n308) );
	nand2_2 U310 ( .x(n193), .a(n268), .b(n267) );
	nand2_5 U311 ( .x(n270), .a(B[29]), .b(A[29]) );
	nand2i_4 U312 ( .x(n328), .a(n102), .b(n162) );
	nand3i_3 U313 ( .x(n329), .a(n290), .b(n328), .c(n320) );
	inv_5 U314 ( .x(n257), .a(n250) );
	mux2i_3 U315 ( .x(n99), .d0(n281), .sl(B[18]), .d1(n278) );
	nand2_3 U316 ( .x(SUM[18]), .a(n99), .b(n100) );
	aoai211_5 U317 ( .x(n133), .a(n239), .b(n240), .c(n57), .d(n270) );
	aoi21_4 U318 ( .x(n129), .a(n130), .b(n131), .c(n132) );
	nand2i_6 U319 ( .x(n231), .a(n77), .b(n232) );
	inv_5 U32 ( .x(n226), .a(B[1]) );
	nor2_8 U320 ( .x(n122), .a(B[19]), .b(A[19]) );
	nor2i_5 U321 ( .x(n297), .a(n55), .b(n183) );
	nor2i_5 U322 ( .x(n296), .a(B[25]), .b(n183) );
	inv_10 U323 ( .x(n233), .a(B[2]) );
	inv_6 U324 ( .x(n232), .a(n227) );
	inv_10 U325 ( .x(n236), .a(B[8]) );
	nand3_4 U326 ( .x(n227), .a(n228), .b(n229), .c(n230) );
	nand2i_4 U327 ( .x(n178), .a(n106), .b(n292) );
	aoai211_3 U328 ( .x(n299), .a(n333), .b(n332), .c(n93), .d(n294) );
	oaoi211_3 U329 ( .x(n93), .a(n96), .b(n95), .c(n321), .d(n94) );
	nor2_2 U33 ( .x(n78), .a(n80), .b(n79) );
	inv_2 U330 ( .x(n311), .a(n77) );
	aoi21_2 U331 ( .x(n77), .a(n310), .b(n81), .c(n78) );
	aoi21_1 U332 ( .x(n340), .a(n197), .b(n342), .c(n341) );
	inv_2 U333 ( .x(n144), .a(n340) );
	inv_0 U334 ( .x(n341), .a(n175) );
	inv_0 U335 ( .x(n342), .a(n256) );
	inv_0 U336 ( .x(n316), .a(n197) );
	nand2_2 U337 ( .x(n256), .a(n73), .b(n257) );
	exnor2_3 U338 ( .x(SUM[29]), .a(n57), .b(n343) );
	inv_2 U339 ( .x(n343), .a(n53) );
	nand2_0 U34 ( .x(n140), .a(B[0]), .b(A[0]) );
	nand2_1 U340 ( .x(n206), .a(n300), .b(n298) );
	mux2i_3 U341 ( .x(SUM[22]), .d0(n280), .sl(n344), .d1(n137) );
	ao21_3 U342 ( .x(n344), .a(n190), .b(n92), .c(n191) );
	inv_2 U343 ( .x(n262), .a(B[13]) );
	aoi21_1 U35 ( .x(n139), .a(n140), .b(n339), .c(n141) );
	nor2i_1 U36 ( .x(n107), .a(n108), .b(n69) );
	inv_2 U37 ( .x(n108), .a(n97) );
	inv_0 U38 ( .x(n103), .a(n254) );
	inv_2 U39 ( .x(n238), .a(A[9]) );
	inv_2 U40 ( .x(n67), .a(B[9]) );
	nand3i_1 U41 ( .x(n320), .a(n289), .b(n254), .c(n162) );
	inv_2 U42 ( .x(n222), .a(A[7]) );
	inv_2 U43 ( .x(n283), .a(n69) );
	ao21_2 U44 ( .x(n199), .a(n200), .b(n283), .c(n97) );
	nor2i_1 U45 ( .x(SUM[0]), .a(n335), .b(n336) );
	inv_2 U46 ( .x(n266), .a(A[11]) );
	nand2i_2 U47 ( .x(n255), .a(B[11]), .b(n266) );
	nor2i_1 U48 ( .x(n151), .a(n152), .b(n153) );
	nand2_1 U49 ( .x(n152), .a(A[14]), .b(B[14]) );
	oaoi211_4 U5 ( .x(n57), .a(A[28]), .b(B[28]), .c(n334), .d(n90) );
	inv_0 U50 ( .x(n153), .a(n252) );
	and2_5 U51 ( .x(n59), .a(n60), .b(n263) );
	inv_4 U52 ( .x(n263), .a(A[14]) );
	nor2i_0 U53 ( .x(n154), .a(n155), .b(n156) );
	nand2_1 U54 ( .x(n155), .a(B[13]), .b(A[13]) );
	inv_5 U55 ( .x(n156), .a(n319) );
	nor2i_0 U56 ( .x(n109), .a(n110), .b(n111) );
	nand2i_2 U57 ( .x(n249), .a(n121), .b(n146) );
	inv_2 U58 ( .x(n259), .a(n249) );
	and2_3 U59 ( .x(n75), .a(n76), .b(n261) );
	aoai211_3 U6 ( .x(n334), .a(n300), .b(n298), .c(n128), .d(n56) );
	inv_0 U60 ( .x(n279), .a(n273) );
	nor2i_0 U61 ( .x(n281), .a(A[18]), .b(n273) );
	nand2i_2 U62 ( .x(n195), .a(A[29]), .b(n240) );
	nor2i_1 U63 ( .x(n170), .a(B[27]), .b(n171) );
	inv_2 U64 ( .x(n171), .a(A[27]) );
	nor2_1 U65 ( .x(n128), .a(B[27]), .b(A[27]) );
	nor2i_1 U66 ( .x(n126), .a(A[26]), .b(n127) );
	inv_2 U67 ( .x(n127), .a(B[26]) );
	inv_2 U68 ( .x(n183), .a(n323) );
	inv_5 U69 ( .x(n98), .a(B[6]) );
	inv_5 U7 ( .x(n72), .a(A[15]) );
	inv_0 U70 ( .x(n66), .a(A[4]) );
	inv_2 U71 ( .x(n285), .a(n105) );
	inv_2 U72 ( .x(n315), .a(n292) );
	nand2i_5 U74 ( .x(n234), .a(n233), .b(n232) );
	exnor2_1 U75 ( .x(SUM[1]), .a(n338), .b(n335) );
	nand2_2 U76 ( .x(n254), .a(n67), .b(n238) );
	inv_2 U77 ( .x(n326), .a(n220) );
	oai21_1 U78 ( .x(n221), .a(n50), .b(n159), .c(n158) );
	inv_2 U79 ( .x(n325), .a(n221) );
	nand2_5 U8 ( .x(n70), .a(n72), .b(n71) );
	nand2_5 U80 ( .x(n319), .a(n68), .b(n262) );
	oai21_1 U81 ( .x(n220), .a(n156), .b(n325), .c(n155) );
	nor2i_1 U82 ( .x(n148), .a(n149), .b(n150) );
	inv_2 U83 ( .x(n150), .a(n146) );
	nand2_1 U84 ( .x(n149), .a(A[16]), .b(B[16]) );
	inv_2 U85 ( .x(n147), .a(n149) );
	nand2i_2 U86 ( .x(n146), .a(B[16]), .b(n260) );
	inv_5 U87 ( .x(n287), .a(n177) );
	nand2i_2 U88 ( .x(n304), .a(A[22]), .b(n116) );
	inv_0 U89 ( .x(n244), .a(A[22]) );
	oai22_1 U90 ( .x(n188), .a(n116), .b(n244), .c(n138), .d(n118) );
	nor2_1 U91 ( .x(n186), .a(n138), .b(n301) );
	inv_2 U92 ( .x(n138), .a(n304) );
	nand2i_0 U93 ( .x(n190), .a(A[21]), .b(n243) );
	inv_0 U94 ( .x(n243), .a(B[21]) );
	inv_0 U95 ( .x(n125), .a(B[24]) );
	nor2i_1 U96 ( .x(n124), .a(A[24]), .b(n125) );
	oai31_2 U97 ( .x(n194), .a(n117), .b(n138), .c(n119), .d(n271) );
	aoi21_1 U98 ( .x(n294), .a(n194), .b(n295), .c(n124) );
	nand2i_2 U99 ( .x(n332), .a(n322), .b(n331) );

endmodule


module EX_DW01_add_32_1_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
	n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
	n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
	n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
	n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
	n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
	n91, n92, n93, n94, n95, n96, n97, n98, n99;


	nor3_1 U10 ( .x(n253), .a(n199), .b(n200), .c(n201) );
	nor3i_1 U100 ( .x(n89), .a(n90), .b(n91), .c(n92) );
	nor2i_1 U102 ( .x(n91), .a(n132), .b(n137) );
	nor3i_1 U103 ( .x(n92), .a(n132), .b(n133), .c(n134) );
	exnor2_1 U104 ( .x(SUM[1]), .a(n82), .b(n249) );
	nand2i_2 U105 ( .x(n218), .a(B[9]), .b(n184) );
	nand2_1 U106 ( .x(n94), .a(A[9]), .b(B[9]) );
	nand3_1 U107 ( .x(n143), .a(n262), .b(n263), .c(n250) );
	nand2i_2 U108 ( .x(n262), .a(n278), .b(n270) );
	nand2i_2 U109 ( .x(n263), .a(n101), .b(n217) );
	inv_2 U11 ( .x(n198), .a(A[24]) );
	nor2_1 U110 ( .x(n250), .a(n135), .b(n181) );
	exor2_1 U111 ( .x(n152), .a(A[15]), .b(B[15]) );
	inv_4 U112 ( .x(n227), .a(n223) );
	nand2i_0 U113 ( .x(n254), .a(n255), .b(n227) );
	inv_0 U114 ( .x(n229), .a(n237) );
	nand2i_0 U115 ( .x(n215), .a(A[14]), .b(n203) );
	inv_2 U116 ( .x(n255), .a(n215) );
	exnor2_1 U117 ( .x(SUM[17]), .a(A[17]), .b(n248) );
	oai21_1 U118 ( .x(n248), .a(n142), .b(n228), .c(A[16]) );
	inv_2 U119 ( .x(n195), .a(A[23]) );
	inv_2 U12 ( .x(n201), .a(A[25]) );
	inv_2 U120 ( .x(n119), .a(n199) );
	nor2i_1 U121 ( .x(n121), .a(A[25]), .b(n199) );
	exor2_1 U122 ( .x(SUM[6]), .a(n75), .b(n98) );
	exnor2_1 U123 ( .x(SUM[12]), .a(n157), .b(n158) );
	exnor2_1 U124 ( .x(SUM[7]), .a(n144), .b(n145) );
	exor2_1 U125 ( .x(SUM[11]), .a(n159), .b(n129) );
	buf_1 U126 ( .x(n54), .a(A[20]) );
	exnor2_1 U127 ( .x(SUM[20]), .a(n54), .b(n247) );
	exnor2_1 U128 ( .x(SUM[14]), .a(n153), .b(n154) );
	exnor2_1 U129 ( .x(SUM[13]), .a(n155), .b(n156) );
	nor2i_0 U13 ( .x(n140), .a(n139), .b(n50) );
	exnor2_1 U130 ( .x(SUM[10]), .a(n160), .b(n161) );
	inv_2 U131 ( .x(n194), .a(A[22]) );
	exnor2_1 U132 ( .x(SUM[22]), .a(n112), .b(n194) );
	exnor2_1 U133 ( .x(SUM[5]), .a(n85), .b(n100) );
	inv_0 U134 ( .x(n188), .a(A[19]) );
	exnor2_1 U135 ( .x(SUM[19]), .a(n108), .b(n188) );
	exor2_1 U136 ( .x(SUM[4]), .a(n70), .b(n103) );
	exnor2_1 U137 ( .x(SUM[8]), .a(n89), .b(n95) );
	exor2_1 U138 ( .x(SUM[9]), .a(n143), .b(n93) );
	exor2_1 U139 ( .x(SUM[15]), .a(n151), .b(n152) );
	inv_4 U14 ( .x(n139), .a(n226) );
	inv_2 U140 ( .x(n200), .a(A[26]) );
	exnor2_1 U141 ( .x(SUM[26]), .a(n120), .b(n200) );
	inv_2 U142 ( .x(n245), .a(A[31]) );
	and2_2 U143 ( .x(n49), .a(n71), .b(n164) );
	inv_6 U145 ( .x(n66), .a(n218) );
	oai21_1 U146 ( .x(n51), .a(n60), .b(n177), .c(n59) );
	inv_1 U148 ( .x(n234), .a(A[28]) );
	exnor2_1 U149 ( .x(SUM[28]), .a(n122), .b(n234) );
	inv_0 U15 ( .x(n202), .a(B[15]) );
	nor2i_1 U150 ( .x(n252), .a(n56), .b(n234) );
	inv_2 U151 ( .x(n55), .a(n234) );
	exnor2_1 U152 ( .x(SUM[29]), .a(n124), .b(n235) );
	inv_2 U153 ( .x(n56), .a(n235) );
	inv_2 U154 ( .x(n235), .a(A[29]) );
	aoi21_1 U155 ( .x(n82), .a(n77), .b(A[1]), .c(n83) );
	and2_2 U156 ( .x(n73), .a(B[1]), .b(A[1]) );
	nand2i_2 U157 ( .x(n258), .a(A[1]), .b(n169) );
	inv_2 U158 ( .x(n57), .a(n128) );
	nand4_1 U159 ( .x(n189), .a(A[19]), .b(A[18]), .c(A[16]), .d(A[17]) );
	nand2i_2 U16 ( .x(n264), .a(A[15]), .b(n202) );
	ao21_1 U160 ( .x(n216), .a(n58), .b(n184), .c(n278) );
	inv_0 U161 ( .x(n58), .a(B[9]) );
	inv_2 U162 ( .x(n184), .a(A[9]) );
	nand2i_2 U163 ( .x(n158), .a(n221), .b(n53) );
	inv_2 U164 ( .x(n221), .a(n267) );
	exor2_1 U165 ( .x(SUM[3]), .a(n146), .b(n147) );
	oai21_2 U166 ( .x(n260), .a(A[3]), .b(n146), .c(B[3]) );
	inv_0 U167 ( .x(n207), .a(A[11]) );
	nand2_0 U168 ( .x(n130), .a(A[11]), .b(B[11]) );
	inv_2 U169 ( .x(n162), .a(A[8]) );
	inv_2 U17 ( .x(n214), .a(n264) );
	nand2_1 U170 ( .x(n186), .a(B[7]), .b(A[7]) );
	inv_2 U171 ( .x(n59), .a(n251) );
	inv_0 U172 ( .x(n60), .a(B[4]) );
	inv_0 U173 ( .x(n180), .a(n177) );
	inv_2 U174 ( .x(n251), .a(n101) );
	inv_2 U175 ( .x(n61), .a(n179) );
	exnor2_1 U176 ( .x(SUM[16]), .a(n149), .b(n150) );
	nand2i_6 U177 ( .x(n149), .a(n138), .b(n78) );
	inv_0 U178 ( .x(n179), .a(B[4]) );
	nor2_0 U179 ( .x(n63), .a(n279), .b(n66) );
	nand2i_2 U18 ( .x(n213), .a(n214), .b(n215) );
	nor2_0 U180 ( .x(n62), .a(n278), .b(n66) );
	nor2_3 U181 ( .x(n65), .a(n136), .b(n66) );
	aoi31_3 U182 ( .x(n72), .a(A[0]), .b(n258), .c(B[0]), .d(n73) );
	nand2_1 U183 ( .x(n99), .a(A[6]), .b(B[6]) );
	inv_5 U184 ( .x(n169), .a(B[1]) );
	inv_2 U185 ( .x(n64), .a(n53) );
	nand2i_1 U186 ( .x(n267), .a(B[12]), .b(n206) );
	inv_0 U187 ( .x(n217), .a(n279) );
	inv_2 U188 ( .x(n128), .a(A[30]) );
	inv_2 U189 ( .x(n67), .a(n238) );
	ao21_1 U19 ( .x(n76), .a(n52), .b(n74), .c(n51) );
	inv_2 U190 ( .x(n68), .a(n224) );
	nand2_0 U191 ( .x(n238), .a(B[13]), .b(A[13]) );
	inv_2 U192 ( .x(n224), .a(n265) );
	inv_0 U193 ( .x(n69), .a(n87) );
	inv_2 U194 ( .x(n70), .a(n69) );
	inv_0 U195 ( .x(n71), .a(B[6]) );
	nand2_0 U196 ( .x(n153), .a(n229), .b(n275) );
	oai221_1 U197 ( .x(n151), .a(n255), .b(n229), .c(n50), .d(n254), .e(n204) );
	nand2_0 U198 ( .x(n249), .a(A[0]), .b(B[0]) );
	exor2_1 U199 ( .x(SUM[0]), .a(A[0]), .b(B[0]) );
	exor2_1 U200 ( .x(n147), .a(B[3]), .b(A[3]) );
	inv_0 U201 ( .x(n83), .a(n258) );
	inv_0 U202 ( .x(n77), .a(n169) );
	aoi211_5 U203 ( .x(n78), .a(n237), .b(n81), .c(n80), .d(n79) );
	inv_2 U204 ( .x(n79), .a(n231) );
	inv_2 U205 ( .x(n81), .a(n213) );
	nand2_0 U206 ( .x(n231), .a(A[15]), .b(B[15]) );
	nand2i_2 U207 ( .x(n230), .a(n204), .b(n264) );
	aoi21_1 U208 ( .x(n90), .a(n251), .b(n132), .c(n182) );
	oai21_2 U209 ( .x(n182), .a(n185), .b(n99), .c(n186) );
	nand2_1 U21 ( .x(n192), .a(n54), .b(A[21]) );
	aoai211_1 U210 ( .x(n159), .a(n268), .b(n269), .c(n211), .d(n209) );
	nand2i_0 U211 ( .x(n161), .a(n211), .b(n209) );
	oai21_1 U212 ( .x(n243), .a(n131), .b(n209), .c(n130) );
	inv_0 U213 ( .x(n203), .a(B[14]) );
	nand2_0 U214 ( .x(n204), .a(A[14]), .b(B[14]) );
	nor2i_0 U215 ( .x(n98), .a(n99), .b(n49) );
	inv_0 U216 ( .x(n261), .a(n99) );
	nand2i_0 U217 ( .x(n265), .a(A[13]), .b(n205) );
	inv_0 U218 ( .x(n205), .a(B[13]) );
	nand2_0 U219 ( .x(n209), .a(B[10]), .b(A[10]) );
	nand2_1 U22 ( .x(n172), .a(B[2]), .b(A[2]) );
	inv_0 U220 ( .x(n208), .a(B[10]) );
	nor2i_5 U221 ( .x(n93), .a(n94), .b(n66) );
	nor2i_3 U222 ( .x(n105), .a(n106), .b(n107) );
	nor2i_3 U223 ( .x(n108), .a(n109), .b(n107) );
	nor2i_3 U224 ( .x(n110), .a(n111), .b(n107) );
	nor2i_3 U225 ( .x(n112), .a(n113), .b(n107) );
	nor2i_3 U226 ( .x(n114), .a(n115), .b(n107) );
	nor2i_3 U227 ( .x(n116), .a(n117), .b(n107) );
	nor2i_3 U228 ( .x(n118), .a(n119), .b(n107) );
	nor2i_3 U229 ( .x(n120), .a(n121), .b(n107) );
	nor2i_1 U23 ( .x(n106), .a(A[17]), .b(n150) );
	nor2i_3 U230 ( .x(n122), .a(n123), .b(n107) );
	nor2i_3 U231 ( .x(n124), .a(n125), .b(n107) );
	nor2_5 U232 ( .x(n126), .a(n127), .b(n128) );
	aoai211_4 U234 ( .x(n146), .a(n171), .b(n170), .c(n72), .d(n172) );
	nand2_5 U235 ( .x(n174), .a(n74), .b(n175) );
	ao21_4 U236 ( .x(n181), .a(n182), .b(n168), .c(n183) );
	inv_6 U237 ( .x(n190), .a(A[21]) );
	nand2i_4 U238 ( .x(n196), .a(n197), .b(n113) );
	nand2i_4 U239 ( .x(n219), .a(n210), .b(n65) );
	nand2i_2 U24 ( .x(n175), .a(n61), .b(n176) );
	nand2i_4 U240 ( .x(n220), .a(n221), .b(n222) );
	nand2i_4 U241 ( .x(n223), .a(n224), .b(n225) );
	nand2i_4 U242 ( .x(n226), .a(n213), .b(n227) );
	exnor2_5 U243 ( .x(SUM[31]), .a(n126), .b(n245) );
	exnor2_5 U244 ( .x(SUM[25]), .a(n118), .b(n201) );
	exnor2_5 U245 ( .x(SUM[24]), .a(n116), .b(n198) );
	exnor2_5 U246 ( .x(SUM[23]), .a(n114), .b(n195) );
	exnor2_5 U247 ( .x(SUM[21]), .a(n110), .b(n190) );
	exnor2_5 U248 ( .x(SUM[18]), .a(n105), .b(n187) );
	nand2_2 U249 ( .x(n197), .a(A[22]), .b(A[23]) );
	inv_2 U25 ( .x(n176), .a(A[4]) );
	nor2i_5 U250 ( .x(n236), .a(n252), .b(n232) );
	nor2i_5 U251 ( .x(n125), .a(n55), .b(n232) );
	nand2i_4 U252 ( .x(n212), .a(B[11]), .b(n207) );
	inv_5 U253 ( .x(n225), .a(n220) );
	inv_5 U254 ( .x(n117), .a(n196) );
	nor2i_5 U255 ( .x(n138), .a(n139), .b(n50) );
	inv_10 U256 ( .x(n107), .a(n149) );
	inv_10 U257 ( .x(n171), .a(B[2]) );
	inv_16 U258 ( .x(n170), .a(A[2]) );
	nand2i_6 U259 ( .x(n127), .a(n107), .b(n236) );
	inv_2 U26 ( .x(n133), .a(n175) );
	nand2i_6 U261 ( .x(n199), .a(n198), .b(n117) );
	inv_7 U263 ( .x(n163), .a(B[7]) );
	nand2i_5 U264 ( .x(n266), .a(A[10]), .b(n208) );
	oai21_1 U265 ( .x(n75), .a(n277), .b(n134), .c(n276) );
	inv_0 U266 ( .x(n276), .a(n51) );
	inv_2 U267 ( .x(n277), .a(n52) );
	or2_1 U268 ( .x(n52), .a(B[4]), .b(A[4]) );
	nand2i_4 U269 ( .x(n134), .a(n102), .b(n87) );
	nand2i_2 U27 ( .x(n232), .a(n233), .b(n119) );
	or2_6 U270 ( .x(n136), .a(n166), .b(n97) );
	or2_1 U271 ( .x(n279), .a(n166), .b(n97) );
	or2_1 U272 ( .x(n278), .a(n166), .b(n97) );
	inv_0 U273 ( .x(n132), .a(n166) );
	nand2i_2 U274 ( .x(n168), .a(B[8]), .b(n162) );
	inv_3 U275 ( .x(n97), .a(n168) );
	nand2i_3 U276 ( .x(n166), .a(n49), .b(n167) );
	nor2_0 U28 ( .x(n135), .a(n279), .b(n137) );
	nand2i_2 U29 ( .x(n137), .a(n179), .b(n180) );
	nor2i_1 U30 ( .x(n142), .a(n139), .b(n50) );
	aoi21_3 U31 ( .x(n50), .a(n52), .b(n74), .c(n51) );
	nor2i_1 U32 ( .x(n111), .a(n54), .b(n189) );
	nor2i_1 U33 ( .x(n115), .a(A[22]), .b(n191) );
	nand2i_2 U34 ( .x(n191), .a(n192), .b(n193) );
	inv_2 U35 ( .x(n113), .a(n191) );
	exor2_1 U36 ( .x(n148), .a(B[2]), .b(A[2]) );
	exnor2_1 U37 ( .x(SUM[2]), .a(n72), .b(n148) );
	inv_0 U38 ( .x(n164), .a(A[6]) );
	inv_5 U40 ( .x(n74), .a(n134) );
	nand2_0 U41 ( .x(n53), .a(A[12]), .b(B[12]) );
	inv_0 U42 ( .x(n206), .a(A[12]) );
	nand2i_0 U43 ( .x(n157), .a(n240), .b(n272) );
	ao21_3 U44 ( .x(n240), .a(n241), .b(n242), .c(n243) );
	nand2i_2 U45 ( .x(n272), .a(n219), .b(n75) );
	nand2i_2 U46 ( .x(n145), .a(n185), .b(n186) );
	inv_2 U47 ( .x(n185), .a(n167) );
	nand2i_3 U48 ( .x(n167), .a(A[7]), .b(n163) );
	nand2i_2 U49 ( .x(n144), .a(n261), .b(n274) );
	nand3_1 U5 ( .x(n233), .a(A[27]), .b(A[26]), .c(A[25]) );
	nand2i_2 U50 ( .x(n274), .a(n49), .b(n76) );
	inv_4 U51 ( .x(n228), .a(n78) );
	oai21_1 U52 ( .x(n246), .a(n140), .b(n228), .c(n253) );
	exnor2_1 U53 ( .x(SUM[27]), .a(A[27]), .b(n246) );
	inv_2 U54 ( .x(n131), .a(n212) );
	nor2i_1 U55 ( .x(n129), .a(n130), .b(n131) );
	inv_0 U56 ( .x(n268), .a(n242) );
	oai21_2 U57 ( .x(n242), .a(n66), .b(n244), .c(n94) );
	inv_2 U58 ( .x(n244), .a(n181) );
	nand2i_2 U59 ( .x(n269), .a(n216), .b(n75) );
	nand2i_2 U6 ( .x(n177), .a(n176), .b(n178) );
	oai21_1 U60 ( .x(n247), .a(n141), .b(n228), .c(n193) );
	nor2i_0 U61 ( .x(n141), .a(n139), .b(n50) );
	inv_2 U62 ( .x(n80), .a(n230) );
	nand2i_2 U63 ( .x(n154), .a(n255), .b(n204) );
	ao21_3 U64 ( .x(n237), .a(n68), .b(n239), .c(n67) );
	nand2i_0 U65 ( .x(n275), .a(n223), .b(n76) );
	nand2i_2 U66 ( .x(n156), .a(n224), .b(n238) );
	nand2i_2 U67 ( .x(n155), .a(n239), .b(n273) );
	ao21_3 U68 ( .x(n239), .a(n267), .b(n240), .c(n64) );
	nand2i_0 U69 ( .x(n273), .a(n220), .b(n76) );
	inv_0 U7 ( .x(n241), .a(n210) );
	inv_2 U70 ( .x(n211), .a(n266) );
	oai211_1 U71 ( .x(n160), .a(n174), .b(n216), .c(n271), .d(n256) );
	nand2i_2 U72 ( .x(n271), .a(n101), .b(n62) );
	aoi21_1 U73 ( .x(n256), .a(n63), .b(n257), .c(n242) );
	inv_2 U74 ( .x(n257), .a(n137) );
	inv_2 U75 ( .x(n270), .a(n174) );
	inv_2 U76 ( .x(n193), .a(n189) );
	nor2i_1 U77 ( .x(n100), .a(n101), .b(n102) );
	nand2_1 U78 ( .x(n101), .a(A[5]), .b(B[5]) );
	inv_2 U79 ( .x(n102), .a(n178) );
	inv_2 U8 ( .x(n222), .a(n219) );
	nand2i_2 U80 ( .x(n178), .a(B[5]), .b(n165) );
	inv_0 U81 ( .x(n165), .a(A[5]) );
	inv_2 U82 ( .x(n173), .a(A[3]) );
	inv_1 U83 ( .x(n259), .a(n146) );
	nand2i_2 U84 ( .x(n86), .a(n61), .b(n176) );
	aoi21_1 U85 ( .x(n85), .a(n86), .b(n70), .c(n88) );
	inv_0 U86 ( .x(n150), .a(A[16]) );
	and3i_1 U87 ( .x(n109), .a(n150), .b(A[18]), .c(A[17]) );
	oai21_2 U88 ( .x(n87), .a(n259), .b(n173), .c(n260) );
	nor2i_1 U89 ( .x(n103), .a(n104), .b(n84) );
	nand2i_2 U9 ( .x(n210), .a(n211), .b(n212) );
	nand2_2 U90 ( .x(n104), .a(n61), .b(A[4]) );
	nor2_1 U91 ( .x(n84), .a(n61), .b(A[4]) );
	inv_2 U92 ( .x(n88), .a(n104) );
	inv_2 U93 ( .x(n187), .a(A[18]) );
	exnor2_3 U94 ( .x(SUM[30]), .a(n127), .b(n57) );
	inv_2 U95 ( .x(n123), .a(n232) );
	inv_2 U96 ( .x(n183), .a(n96) );
	nand2_0 U98 ( .x(n96), .a(A[8]), .b(B[8]) );
	nor2i_1 U99 ( .x(n95), .a(n96), .b(n97) );

endmodule


module EX_DW01_cmp2_32_3_test_1 (  A, B, LEQ, TC, LT_LE, GE_GT );

input  LEQ, TC;
input [31:0] A, B;
output  LT_LE, GE_GT;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n15, n16,
	n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
	n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
	n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
	n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
	n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
	n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	nand2i_2 U10 ( .x(n76), .a(n107), .b(n123) );
	inv_2 U100 ( .x(n72), .a(A[28]) );
	oa22_1 U101 ( .x(n15), .a(B[15]), .b(n62), .c(B[16]), .d(n61) );
	oai22_1 U102 ( .x(n37), .a(A[14]), .b(n64), .c(A[15]), .d(n63) );
	nand2i_2 U105 ( .x(n137), .a(A[24]), .b(B[24]) );
	inv_2 U106 ( .x(n17), .a(n49) );
	inv_2 U107 ( .x(n49), .a(A[1]) );
	inv_2 U108 ( .x(n19), .a(n18) );
	inv_2 U109 ( .x(n18), .a(B[30]) );
	inv_2 U110 ( .x(n66), .a(B[19]) );
	nand4_1 U111 ( .x(n71), .a(A[17]), .b(n102), .c(n101), .d(n65) );
	aoi22_1 U112 ( .x(n124), .a(A[30]), .b(n18), .c(A[29]), .d(n73) );
	oai22_1 U114 ( .x(n142), .a(B[6]), .b(n94), .c(B[5]), .d(n93) );
	aoi21_1 U115 ( .x(n68), .a(A[20]), .b(n26), .c(n106) );
	aoi22_1 U116 ( .x(n119), .a(A[13]), .b(n53), .c(A[14]), .d(n64) );
	inv_1 U117 ( .x(n56), .a(B[8]) );
	nor2i_0 U118 ( .x(n27), .a(A[8]), .b(B[8]) );
	inv_0 U119 ( .x(n91), .a(A[11]) );
	nor2i_0 U120 ( .x(n34), .a(B[11]), .b(A[11]) );
	nor2i_0 U121 ( .x(n33), .a(B[3]), .b(A[3]) );
	inv_0 U122 ( .x(n97), .a(A[0]) );
	inv_0 U123 ( .x(n129), .a(B[7]) );
	oai22_1 U124 ( .x(n117), .a(B[7]), .b(n136), .c(n136), .d(n48) );
	inv_0 U125 ( .x(n55), .a(A[9]) );
	oai22_1 U126 ( .x(n143), .a(A[9]), .b(n57), .c(A[8]), .d(n56) );
	inv_0 U127 ( .x(n53), .a(B[13]) );
	and3i_3 U128 ( .x(LT_LE), .a(n22), .b(n20), .c(n21) );
	nand3_3 U129 ( .x(n74), .a(n75), .b(n76), .c(n77) );
	nand2i_3 U13 ( .x(n121), .a(B[27]), .b(A[27]) );
	nand4_1 U130 ( .x(n38), .a(n101), .b(n102), .c(n103), .d(n104) );
	nor3i_5 U131 ( .x(n79), .a(n115), .b(n112), .c(n74) );
	aoi22_3 U132 ( .x(n21), .a(n130), .b(n131), .c(n96), .d(n130) );
	aoi22_3 U133 ( .x(n20), .a(n132), .b(n130), .c(n133), .d(n130) );
	nand4_1 U134 ( .x(n46), .a(A[23]), .b(n114), .c(n137), .d(n60) );
	nand4_1 U135 ( .x(n144), .a(n145), .b(n15), .c(n119), .d(n139) );
	nand2i_5 U136 ( .x(n69), .a(B[22]), .b(A[22]) );
	nand2i_5 U137 ( .x(n107), .a(A[27]), .b(B[27]) );
	inv_0 U138 ( .x(n89), .a(A[29]) );
	nand3i_2 U139 ( .x(n22), .a(n39), .b(n134), .c(n135) );
	nand3_1 U14 ( .x(n75), .a(n121), .b(n108), .c(n123) );
	inv_0 U140 ( .x(n62), .a(A[15]) );
	nand2i_1 U141 ( .x(n141), .a(A[6]), .b(B[6]) );
	inv_0 U142 ( .x(n92), .a(A[23]) );
	nand2i_4 U143 ( .x(n123), .a(B[28]), .b(A[28]) );
	nor2i_2 U144 ( .x(n108), .a(B[26]), .b(A[26]) );
	nor2i_0 U145 ( .x(n120), .a(A[24]), .b(B[24]) );
	nand2i_2 U15 ( .x(n114), .a(A[25]), .b(B[25]) );
	nor2i_1 U16 ( .x(n100), .a(n19), .b(A[30]) );
	nand2i_0 U17 ( .x(n24), .a(A[20]), .b(n99) );
	nand2i_2 U18 ( .x(n98), .a(A[21]), .b(B[21]) );
	nor2i_1 U19 ( .x(n105), .a(A[18]), .b(B[18]) );
	nand2i_2 U20 ( .x(n99), .a(B[21]), .b(A[21]) );
	nand2i_2 U21 ( .x(n104), .a(A[16]), .b(B[16]) );
	nand2i_0 U22 ( .x(n103), .a(A[17]), .b(B[17]) );
	nand2i_2 U23 ( .x(n102), .a(A[18]), .b(B[18]) );
	nand2i_2 U24 ( .x(n101), .a(A[19]), .b(B[19]) );
	nand2i_2 U25 ( .x(n113), .a(A[31]), .b(B[31]) );
	nand2i_2 U26 ( .x(n126), .a(B[31]), .b(A[31]) );
	inv_2 U27 ( .x(n73), .a(B[29]) );
	nand3_1 U28 ( .x(n47), .a(n121), .b(n122), .c(n123) );
	inv_2 U29 ( .x(n60), .a(B[23]) );
	aoi21_1 U30 ( .x(n45), .a(n120), .b(n114), .c(n35) );
	and3i_1 U31 ( .x(n44), .a(n47), .b(n45), .c(n46) );
	inv_0 U32 ( .x(n90), .a(A[12]) );
	oai22_1 U33 ( .x(n138), .a(B[11]), .b(n91), .c(B[12]), .d(n90) );
	nand2_2 U34 ( .x(n139), .a(n16), .b(n138) );
	and3i_1 U35 ( .x(n28), .a(n31), .b(n29), .c(n30) );
	nand2i_0 U36 ( .x(n29), .a(B[3]), .b(A[3]) );
	nand2i_2 U37 ( .x(n30), .a(B[2]), .b(A[2]) );
	nand3_1 U38 ( .x(n31), .a(n87), .b(n97), .c(n88) );
	oai211_1 U39 ( .x(n118), .a(n32), .b(n33), .c(n29), .d(n87) );
	nor2i_0 U40 ( .x(n32), .a(B[2]), .b(A[2]) );
	nand2i_2 U41 ( .x(n87), .a(B[4]), .b(A[4]) );
	inv_2 U42 ( .x(n136), .a(n141) );
	or3i_2 U43 ( .x(n116), .a(n95), .b(n132), .c(n133) );
	and3i_1 U44 ( .x(n95), .a(n96), .b(n49), .c(B[1]) );
	nand2i_0 U45 ( .x(n81), .a(A[10]), .b(B[10]) );
	oa22_1 U46 ( .x(n16), .a(A[13]), .b(n53), .c(A[12]), .d(n52) );
	inv_2 U47 ( .x(n52), .a(B[12]) );
	nand2_2 U48 ( .x(n80), .a(n140), .b(n143) );
	inv_2 U49 ( .x(n140), .a(n58) );
	oai22_1 U50 ( .x(n58), .a(B[9]), .b(n55), .c(B[10]), .d(n54) );
	inv_2 U51 ( .x(n57), .a(B[9]) );
	nand2_2 U52 ( .x(n112), .a(n113), .b(n114) );
	nand2_2 U53 ( .x(n115), .a(n100), .b(n126) );
	inv_0 U54 ( .x(n26), .a(B[20]) );
	nor3_1 U55 ( .x(n23), .a(n24), .b(n25), .c(n26) );
	inv_0 U56 ( .x(n59), .a(B[22]) );
	oai22_1 U57 ( .x(n109), .a(A[22]), .b(n59), .c(n25), .d(n98) );
	inv_2 U58 ( .x(n111), .a(n137) );
	aoi21_1 U59 ( .x(n110), .a(B[23]), .b(n92), .c(n111) );
	nand2i_2 U6 ( .x(n122), .a(B[26]), .b(A[26]) );
	nor3i_1 U60 ( .x(n78), .a(n110), .b(n109), .c(n23) );
	inv_2 U61 ( .x(n25), .a(n69) );
	inv_0 U62 ( .x(n65), .a(B[17]) );
	aoi22_1 U63 ( .x(n70), .a(A[19]), .b(n66), .c(n105), .d(n101) );
	inv_2 U64 ( .x(n106), .a(n99) );
	nand4_1 U65 ( .x(n67), .a(n68), .b(n69), .c(n70), .d(n71) );
	inv_0 U66 ( .x(n63), .a(B[15]) );
	inv_2 U67 ( .x(n64), .a(B[14]) );
	aoi21_1 U68 ( .x(n36), .a(n15), .b(n37), .c(n38) );
	nand2i_2 U69 ( .x(n135), .a(n88), .b(n130) );
	nor2i_1 U7 ( .x(n35), .a(A[25]), .b(B[25]) );
	nand2i_2 U70 ( .x(n88), .a(B[1]), .b(n17) );
	inv_2 U71 ( .x(n84), .a(n43) );
	aoai211_1 U72 ( .x(n134), .a(n84), .b(n144), .c(n125), .d(n127) );
	inv_2 U73 ( .x(n145), .a(n67) );
	oai211_1 U74 ( .x(n125), .a(n44), .b(n74), .c(n124), .d(n126) );
	nor2i_1 U75 ( .x(n127), .a(n115), .b(n128) );
	inv_2 U76 ( .x(n128), .a(n113) );
	aoi211_1 U77 ( .x(n39), .a(n40), .b(n41), .c(n42), .d(n43) );
	nand2_2 U78 ( .x(n40), .a(n142), .b(n117) );
	aoi211_1 U79 ( .x(n41), .a(A[7]), .b(n129), .c(n27), .d(n58) );
	oai211_3 U80 ( .x(n43), .a(n36), .b(n67), .c(n78), .d(n79) );
	inv_5 U81 ( .x(n130), .a(n82) );
	and4i_1 U82 ( .x(n86), .a(n28), .b(n116), .c(n117), .d(n118) );
	nand4i_1 U83 ( .x(n42), .a(n34), .b(n80), .c(n16), .d(n81) );
	inv_2 U84 ( .x(n85), .a(n42) );
	inv_2 U85 ( .x(n50), .a(B[4]) );
	inv_2 U86 ( .x(n51), .a(B[5]) );
	oai22_1 U87 ( .x(n83), .a(A[5]), .b(n51), .c(A[4]), .d(n50) );
	nand4i_1 U88 ( .x(n82), .a(n83), .b(n84), .c(n85), .d(n86) );
	inv_0 U89 ( .x(n54), .a(A[10]) );
	aoi22_1 U9 ( .x(n77), .a(B[29]), .b(n89), .c(B[28]), .d(n72) );
	inv_2 U90 ( .x(n132), .a(n29) );
	inv_2 U91 ( .x(n133), .a(n30) );
	inv_2 U92 ( .x(n131), .a(B[0]) );
	inv_2 U93 ( .x(n96), .a(n87) );
	inv_0 U95 ( .x(n61), .a(A[16]) );
	inv_0 U96 ( .x(n93), .a(A[5]) );
	inv_2 U97 ( .x(n48), .a(A[7]) );
	inv_0 U99 ( .x(n94), .a(A[6]) );

endmodule


module EX_DW01_cmp2_32_0 (  A, B, LEQ, TC, LT_LE, GE_GT );

input  LEQ, TC;
input [31:0] A, B;
output  LT_LE, GE_GT;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n15, n150, n151, n152, n153, n154, n155, n156, n157, n158,
	n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
	n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
	n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57,
	n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
	n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
	n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	aoi211_1 U10 ( .x(n81), .a(A[20]), .b(n62), .c(n110), .d(n112) );
	oa22_2 U100 ( .x(n16), .a(A[31]), .b(n54), .c(A[30]), .d(n53) );
	nand2_2 U101 ( .x(n45), .a(n17), .b(B[11]) );
	inv_0 U102 ( .x(n17), .a(A[11]) );
	inv_2 U103 ( .x(n18), .a(n62) );
	inv_2 U104 ( .x(n62), .a(B[20]) );
	inv_2 U105 ( .x(n84), .a(A[3]) );
	inv_2 U106 ( .x(n19), .a(n53) );
	inv_2 U107 ( .x(n53), .a(B[30]) );
	inv_2 U108 ( .x(n21), .a(n20) );
	inv_0 U109 ( .x(n65), .a(B[13]) );
	nand2i_2 U11 ( .x(n131), .a(B[22]), .b(A[22]) );
	inv_0 U110 ( .x(n22), .a(n75) );
	inv_2 U111 ( .x(n76), .a(n68) );
	nand2_2 U112 ( .x(n75), .a(n99), .b(n100) );
	inv_2 U113 ( .x(n74), .a(n45) );
	oai22_1 U114 ( .x(n27), .a(B[5]), .b(n28), .c(B[6]), .d(n25) );
	nand4_1 U115 ( .x(n82), .a(A[17]), .b(n97), .c(n98), .d(n94) );
	nor2i_0 U116 ( .x(n128), .a(B[17]), .b(A[17]) );
	inv_0 U117 ( .x(n28), .a(A[5]) );
	nand2i_0 U118 ( .x(n127), .a(A[5]), .b(B[5]) );
	inv_1 U119 ( .x(n71), .a(B[8]) );
	aoi22_1 U12 ( .x(n80), .a(A[19]), .b(n78), .c(n116), .d(n98) );
	inv_0 U120 ( .x(n92), .a(B[3]) );
	nand2i_0 U121 ( .x(n107), .a(B[24]), .b(A[24]) );
	oai22_1 U122 ( .x(n60), .a(A[25]), .b(n56), .c(A[24]), .d(n55) );
	oai31_1 U123 ( .x(n132), .a(n42), .b(n118), .c(n133), .d(n130) );
	oai222_1 U124 ( .x(n134), .a(n42), .b(n126), .c(n42), .d(n120), .e(n42),
		.f(n122) );
	oai31_1 U125 ( .x(n138), .a(n42), .b(n127), .c(n27), .d(n135) );
	oai21_1 U126 ( .x(n142), .a(n24), .b(n42), .c(n143) );
	nor2_2 U127 ( .x(n41), .a(n42), .b(n43) );
	oai21_1 U128 ( .x(n146), .a(n42), .b(n77), .c(n147) );
	aoi22_1 U129 ( .x(n24), .a(B[6]), .b(n25), .c(B[7]), .d(n26) );
	inv_2 U13 ( .x(n78), .a(B[19]) );
	nand2i_0 U130 ( .x(n113), .a(B[7]), .b(A[7]) );
	nand2i_0 U131 ( .x(n114), .a(B[8]), .b(A[8]) );
	oai22_1 U132 ( .x(n100), .a(A[9]), .b(n72), .c(A[8]), .d(n71) );
	nand4i_1 U133 ( .x(n73), .a(n74), .b(n75), .c(n76), .d(n77) );
	inv_2 U134 ( .x(n115), .a(n77) );
	nand2i_4 U135 ( .x(n77), .a(A[10]), .b(B[10]) );
	nor2i_0 U136 ( .x(n108), .a(B[21]), .b(A[21]) );
	inv_0 U137 ( .x(n63), .a(A[16]) );
	nand2i_0 U138 ( .x(n129), .a(A[16]), .b(B[16]) );
	inv_0 U139 ( .x(n31), .a(A[14]) );
	nor2i_1 U14 ( .x(n116), .a(A[18]), .b(B[18]) );
	aoi222_1 U140 ( .x(n90), .a(n76), .b(n117), .c(A[13]), .d(n65), .e(A[14]),
		.f(n93) );
	inv_0 U141 ( .x(n66), .a(A[12]) );
	oai22_1 U142 ( .x(n68), .a(A[13]), .b(n65), .c(A[12]), .d(n64) );
	inv_0 U143 ( .x(n25), .a(A[6]) );
	inv_0 U144 ( .x(n70), .a(A[10]) );
	aoi21_3 U145 ( .x(LT_LE), .a(n50), .b(n51), .c(n52) );
	nor3i_5 U146 ( .x(n89), .a(n15), .b(n44), .c(n33) );
	nand2i_4 U147 ( .x(n144), .a(n142), .b(n141) );
	nor3_4 U148 ( .x(n50), .a(n144), .b(n145), .c(n146) );
	nand4_5 U149 ( .x(n42), .a(n88), .b(n89), .c(n90), .d(n91) );
	nand2i_0 U15 ( .x(n158), .a(B[21]), .b(A[21]) );
	nand3i_5 U150 ( .x(n120), .a(A[0]), .b(n119), .c(n121) );
	oai22_1 U16 ( .x(n86), .a(B[3]), .b(n84), .c(B[4]), .d(n83) );
	nand2i_2 U17 ( .x(n157), .a(B[1]), .b(A[1]) );
	or3i_2 U18 ( .x(n155), .a(n123), .b(n156), .c(A[2]) );
	aoi21_1 U19 ( .x(n58), .a(n104), .b(n101), .c(n39) );
	nor2i_1 U20 ( .x(n104), .a(n21), .b(A[27]) );
	nor2i_1 U21 ( .x(n39), .a(B[28]), .b(A[28]) );
	nand3_1 U22 ( .x(n57), .a(n49), .b(n105), .c(n101) );
	inv_0 U23 ( .x(n20), .a(B[27]) );
	nor2i_1 U24 ( .x(n105), .a(B[26]), .b(A[26]) );
	nor2i_1 U25 ( .x(n40), .a(B[29]), .b(A[29]) );
	nand2i_2 U26 ( .x(n140), .a(A[23]), .b(B[23]) );
	nand2i_2 U27 ( .x(n97), .a(A[18]), .b(B[18]) );
	oai31_2 U28 ( .x(n121), .a(n87), .b(n156), .c(n86), .d(n155) );
	inv_2 U29 ( .x(n96), .a(B[0]) );
	nand3i_1 U30 ( .x(n43), .a(n96), .b(n119), .c(n121) );
	nand2i_2 U31 ( .x(n98), .a(A[19]), .b(B[19]) );
	nand2i_2 U32 ( .x(n91), .a(n113), .b(n154) );
	inv_2 U33 ( .x(n154), .a(n73) );
	inv_2 U34 ( .x(n93), .a(B[14]) );
	inv_0 U35 ( .x(n67), .a(A[11]) );
	oai22_1 U36 ( .x(n117), .a(B[11]), .b(n67), .c(B[12]), .d(n66) );
	nand3_1 U37 ( .x(n33), .a(n80), .b(n81), .c(n82) );
	and3i_1 U38 ( .x(n44), .a(n47), .b(n45), .c(n46) );
	nand2i_2 U39 ( .x(n88), .a(n114), .b(n154) );
	nor2_1 U40 ( .x(n37), .a(n35), .b(n38) );
	nand2i_2 U41 ( .x(n38), .a(B[26]), .b(A[26]) );
	nor2_1 U42 ( .x(n34), .a(n35), .b(n36) );
	nand2i_2 U43 ( .x(n36), .a(B[25]), .b(A[25]) );
	nand2i_2 U44 ( .x(n152), .a(B[31]), .b(A[31]) );
	nand2i_2 U45 ( .x(n101), .a(B[28]), .b(A[28]) );
	nor2_1 U46 ( .x(n48), .a(n35), .b(n49) );
	nand4i_1 U47 ( .x(n35), .a(n40), .b(n57), .c(n58), .d(n16) );
	nand2i_2 U48 ( .x(n49), .a(n21), .b(A[27]) );
	nor2i_1 U49 ( .x(n103), .a(A[29]), .b(B[29]) );
	inv_2 U50 ( .x(n54), .a(B[31]) );
	nor2i_1 U51 ( .x(n102), .a(A[30]), .b(n19) );
	nor2i_1 U52 ( .x(n106), .a(A[23]), .b(B[23]) );
	aoi211_1 U53 ( .x(n135), .a(n128), .b(n136), .c(n137), .d(n32) );
	oai22_1 U54 ( .x(n137), .a(A[22]), .b(n95), .c(n33), .d(n129) );
	inv_0 U55 ( .x(n95), .a(B[22]) );
	nor3i_1 U56 ( .x(n32), .a(n15), .b(n29), .c(n33) );
	aoi22_1 U57 ( .x(n130), .a(n108), .b(n131), .c(n111), .d(n109) );
	nor2i_1 U58 ( .x(n111), .a(n18), .b(n112) );
	inv_2 U59 ( .x(n112), .a(n158) );
	nand2i_2 U6 ( .x(n47), .a(n115), .b(n76) );
	nor2i_1 U60 ( .x(n109), .a(n79), .b(n110) );
	inv_0 U61 ( .x(n79), .a(A[20]) );
	inv_2 U62 ( .x(n110), .a(n131) );
	inv_2 U63 ( .x(n85), .a(A[1]) );
	nand3_1 U64 ( .x(n118), .a(n119), .b(n85), .c(B[1]) );
	oai22_1 U65 ( .x(n124), .a(A[3]), .b(n92), .c(A[2]), .d(n87) );
	inv_2 U66 ( .x(n119), .a(n27) );
	inv_2 U67 ( .x(n83), .a(A[4]) );
	inv_2 U68 ( .x(n123), .a(n86) );
	nand3_1 U69 ( .x(n122), .a(n123), .b(n119), .c(n124) );
	inv_0 U7 ( .x(n30), .a(A[15]) );
	inv_2 U70 ( .x(n156), .a(n157) );
	inv_2 U71 ( .x(n87), .a(B[2]) );
	nand2i_2 U72 ( .x(n125), .a(A[4]), .b(B[4]) );
	nand2i_2 U73 ( .x(n126), .a(n125), .b(n119) );
	nand2i_2 U74 ( .x(n59), .a(n60), .b(n61) );
	inv_2 U75 ( .x(n56), .a(B[25]) );
	inv_2 U76 ( .x(n55), .a(B[24]) );
	inv_2 U77 ( .x(n72), .a(B[9]) );
	inv_0 U78 ( .x(n69), .a(A[9]) );
	oai22_1 U79 ( .x(n46), .a(B[10]), .b(n70), .c(B[9]), .d(n69) );
	aoi22_1 U8 ( .x(n29), .a(B[15]), .b(n30), .c(B[14]), .d(n31) );
	inv_4 U80 ( .x(n99), .a(n46) );
	inv_2 U81 ( .x(n64), .a(B[12]) );
	nor2_1 U82 ( .x(n141), .a(n41), .b(n139) );
	oai21_1 U83 ( .x(n139), .a(n33), .b(n97), .c(n140) );
	inv_0 U84 ( .x(n26), .a(A[7]) );
	nand2i_2 U85 ( .x(n143), .a(n98), .b(n136) );
	inv_2 U86 ( .x(n136), .a(n33) );
	nand4_1 U87 ( .x(n52), .a(n148), .b(n149), .c(n150), .d(n151) );
	aoi222_1 U88 ( .x(n148), .a(n106), .b(n147), .c(n102), .d(n16), .e(n103),
		.f(n16) );
	nand2i_2 U89 ( .x(n149), .a(n107), .b(n147) );
	inv_2 U9 ( .x(n94), .a(B[17]) );
	aoi21_1 U90 ( .x(n150), .a(n153), .b(n61), .c(n48) );
	inv_2 U91 ( .x(n153), .a(n101) );
	inv_2 U92 ( .x(n61), .a(n35) );
	nor3i_1 U93 ( .x(n151), .a(n152), .b(n34), .c(n37) );
	nor3_1 U94 ( .x(n51), .a(n134), .b(n132), .c(n138) );
	inv_2 U95 ( .x(n133), .a(n121) );
	inv_2 U96 ( .x(n147), .a(n59) );
	inv_5 U97 ( .x(n23), .a(n42) );
	ao222_2 U98 ( .x(n145), .a(n23), .b(n22), .c(n68), .d(n23), .e(n23), .f(n74) );
	oa22_1 U99 ( .x(n15), .a(B[15]), .b(n30), .c(B[16]), .d(n63) );

endmodule


module EX_DW01_cmp2_32_5_test_1 (  A, B, LEQ, TC, LT_LE, GE_GT );

input  LEQ, TC;
input [31:0] A, B;
output  LT_LE, GE_GT;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n15, n16, n17, n18, n19, n20, n21,
	n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
	n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
	n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
	n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
	n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
	n92, n93, n94, n95, n96, n97, n98, n99;


	nand3_1 U10 ( .x(n75), .a(n136), .b(n105), .c(n137) );
	inv_2 U100 ( .x(n21), .a(n88) );
	inv_2 U101 ( .x(n22), .a(A[28]) );
	aoi22_1 U102 ( .x(n67), .a(A[19]), .b(n65), .c(n103), .d(n99) );
	nand4i_4 U103 ( .x(n42), .a(n19), .b(n66), .c(n67), .d(n68) );
	inv_0 U104 ( .x(n64), .a(B[17]) );
	nand2_0 U105 ( .x(n86), .a(n24), .b(A[3]) );
	oai22_1 U106 ( .x(n123), .a(B[30]), .b(n88), .c(B[29]), .d(n89) );
	inv_0 U107 ( .x(n94), .a(A[6]) );
	inv_0 U108 ( .x(n58), .a(B[20]) );
	oai22_1 U109 ( .x(n140), .a(A[9]), .b(n57), .c(A[8]), .d(n56) );
	nor2i_0 U110 ( .x(n31), .a(A[8]), .b(B[8]) );
	aoi22_1 U111 ( .x(n26), .a(A[0]), .b(n128), .c(n129), .d(n128) );
	nand2i_2 U112 ( .x(n66), .a(B[22]), .b(A[22]) );
	oai22_1 U113 ( .x(n139), .a(B[11]), .b(n91), .c(B[12]), .d(n90) );
	nor2i_0 U114 ( .x(n34), .a(B[11]), .b(A[11]) );
	nor2i_0 U115 ( .x(n33), .a(B[3]), .b(A[3]) );
	inv_0 U116 ( .x(n131), .a(B[0]) );
	aoi221_1 U117 ( .x(n47), .a(n18), .b(n48), .c(A[7]), .d(n49), .e(n50) );
	nand2i_2 U118 ( .x(n100), .a(A[18]), .b(B[18]) );
	inv_0 U119 ( .x(n57), .a(B[9]) );
	inv_2 U12 ( .x(n122), .a(n136) );
	aoi22_1 U120 ( .x(n40), .a(A[13]), .b(n53), .c(A[14]), .d(n63) );
	and3i_3 U121 ( .x(LT_LE), .a(n27), .b(n25), .c(n26) );
	aoi21_3 U122 ( .x(n36), .a(n15), .b(n37), .c(n38) );
	oai211_4 U123 ( .x(n44), .a(n36), .b(n42), .c(n76), .d(n77) );
	nand4i_4 U124 ( .x(n81), .a(n82), .b(n83), .c(n18), .d(n84) );
	nor2i_5 U125 ( .x(n96), .a(B[21]), .b(A[21]) );
	nand4_1 U126 ( .x(n38), .a(n99), .b(n100), .c(n101), .d(n102) );
	nand2i_4 U127 ( .x(n106), .a(A[27]), .b(B[27]) );
	and4i_5 U128 ( .x(n77), .a(n72), .b(n110), .c(n111), .d(n112) );
	nand4_1 U129 ( .x(n82), .a(n113), .b(n114), .c(n115), .d(n116) );
	nand2i_2 U13 ( .x(n74), .a(n106), .b(n137) );
	nand2i_4 U130 ( .x(n97), .a(B[21]), .b(A[21]) );
	nand4_1 U131 ( .x(n113), .a(n95), .b(n85), .c(n86), .d(n87) );
	inv_10 U132 ( .x(n61), .a(A[15]) );
	nand2i_6 U133 ( .x(n136), .a(B[27]), .b(A[27]) );
	inv_3 U134 ( .x(n70), .a(B[28]) );
	nand2i_1 U135 ( .x(n137), .a(B[28]), .b(n23) );
	nor2i_0 U136 ( .x(n105), .a(B[26]), .b(A[26]) );
	nand2i_0 U137 ( .x(n110), .a(A[24]), .b(B[24]) );
	oai22_1 U15 ( .x(n73), .a(A[29]), .b(n71), .c(n23), .d(n70) );
	inv_0 U16 ( .x(n71), .a(B[29]) );
	inv_2 U17 ( .x(n23), .a(n22) );
	inv_2 U18 ( .x(n90), .a(A[12]) );
	inv_2 U19 ( .x(n91), .a(A[11]) );
	inv_2 U20 ( .x(n55), .a(A[9]) );
	inv_2 U21 ( .x(n54), .a(A[10]) );
	nand2i_1 U22 ( .x(n29), .a(n58), .b(n97) );
	nor3_1 U23 ( .x(n28), .a(n29), .b(A[20]), .c(n30) );
	nand2i_2 U24 ( .x(n120), .a(A[25]), .b(B[25]) );
	inv_2 U25 ( .x(n109), .a(n120) );
	inv_2 U26 ( .x(n92), .a(A[23]) );
	aoi21_1 U27 ( .x(n108), .a(B[23]), .b(n92), .c(n109) );
	aoi21_1 U28 ( .x(n107), .a(n96), .b(n66), .c(n35) );
	nor2i_0 U29 ( .x(n35), .a(B[22]), .b(A[22]) );
	nand4_1 U30 ( .x(n68), .a(n100), .b(n64), .c(n99), .d(A[17]) );
	nor2i_1 U31 ( .x(n103), .a(A[18]), .b(B[18]) );
	inv_2 U32 ( .x(n30), .a(n66) );
	inv_2 U33 ( .x(n104), .a(n97) );
	nand2i_0 U34 ( .x(n102), .a(A[16]), .b(B[16]) );
	nand2i_0 U35 ( .x(n101), .a(A[17]), .b(B[17]) );
	nand2i_2 U36 ( .x(n99), .a(A[19]), .b(B[19]) );
	oai22_1 U37 ( .x(n37), .a(A[14]), .b(n63), .c(A[15]), .d(n62) );
	nor2i_0 U38 ( .x(n32), .a(B[2]), .b(A[2]) );
	nor2i_1 U39 ( .x(n95), .a(n20), .b(A[1]) );
	inv_0 U40 ( .x(n69), .a(B[26]) );
	nand2i_0 U41 ( .x(n87), .a(B[2]), .b(A[2]) );
	nand2i_0 U42 ( .x(n117), .a(n20), .b(A[1]) );
	nand2i_2 U43 ( .x(n50), .a(n31), .b(n17) );
	inv_0 U44 ( .x(n93), .a(A[5]) );
	oai22_1 U45 ( .x(n48), .a(B[6]), .b(n94), .c(B[5]), .d(n93) );
	nand2_2 U46 ( .x(n112), .a(n98), .b(n135) );
	nand2i_2 U47 ( .x(n111), .a(A[31]), .b(B[31]) );
	inv_2 U48 ( .x(n127), .a(n111) );
	nand2i_2 U49 ( .x(n46), .a(n127), .b(n112) );
	inv_2 U50 ( .x(n89), .a(A[29]) );
	inv_2 U51 ( .x(n88), .a(A[30]) );
	nand2i_2 U52 ( .x(n135), .a(B[31]), .b(A[31]) );
	inv_2 U53 ( .x(n126), .a(n135) );
	inv_2 U54 ( .x(n141), .a(n137) );
	nand4i_1 U55 ( .x(n125), .a(n141), .b(n121), .c(n119), .d(n138) );
	nand3i_1 U56 ( .x(n72), .a(n73), .b(n74), .c(n75) );
	inv_2 U57 ( .x(n124), .a(n72) );
	aoi211_1 U58 ( .x(n45), .a(n124), .b(n125), .c(n126), .d(n123) );
	nand2_0 U59 ( .x(n41), .a(n16), .b(n139) );
	nor2i_0 U6 ( .x(n98), .a(B[30]), .b(n21) );
	inv_2 U60 ( .x(n60), .a(A[16]) );
	oa22_1 U61 ( .x(n15), .a(B[15]), .b(n61), .c(B[16]), .d(n60) );
	and4i_1 U62 ( .x(n39), .a(n42), .b(n15), .c(n40), .d(n41) );
	inv_2 U63 ( .x(n84), .a(n78) );
	nand2i_0 U64 ( .x(n80), .a(A[10]), .b(B[10]) );
	inv_0 U65 ( .x(n52), .a(B[12]) );
	nand2_2 U66 ( .x(n79), .a(n17), .b(n140) );
	nand4i_1 U67 ( .x(n78), .a(n34), .b(n79), .c(n16), .d(n80) );
	and3i_1 U68 ( .x(n76), .a(n28), .b(n107), .c(n108) );
	inv_5 U69 ( .x(n83), .a(n44) );
	nand4i_1 U7 ( .x(n138), .a(B[23]), .b(n120), .c(A[23]), .d(n110) );
	oai211_1 U70 ( .x(n116), .a(n32), .b(n33), .c(n86), .d(n85) );
	nand2i_0 U71 ( .x(n115), .a(A[4]), .b(B[4]) );
	nand2i_0 U72 ( .x(n114), .a(A[5]), .b(B[5]) );
	nand4i_1 U73 ( .x(n27), .a(n43), .b(n132), .c(n133), .d(n134) );
	oaoi211_1 U74 ( .x(n43), .a(n39), .b(n44), .c(n45), .d(n46) );
	or3i_2 U75 ( .x(n132), .a(n83), .b(n78), .c(n47) );
	nand2i_2 U76 ( .x(n133), .a(n117), .b(n128) );
	inv_5 U77 ( .x(n128), .a(n81) );
	nand2i_2 U78 ( .x(n134), .a(n87), .b(n128) );
	inv_2 U79 ( .x(n129), .a(n85) );
	aoi22_1 U8 ( .x(n119), .a(A[25]), .b(n59), .c(n118), .d(n120) );
	nand2i_2 U80 ( .x(n85), .a(B[4]), .b(A[4]) );
	aoi22_1 U81 ( .x(n25), .a(n130), .b(n128), .c(n128), .d(n131) );
	inv_2 U82 ( .x(n130), .a(n86) );
	inv_0 U83 ( .x(n53), .a(B[13]) );
	inv_2 U84 ( .x(n59), .a(B[25]) );
	inv_2 U85 ( .x(n49), .a(B[7]) );
	inv_0 U86 ( .x(n65), .a(B[19]) );
	inv_0 U87 ( .x(n63), .a(B[14]) );
	inv_0 U88 ( .x(n56), .a(B[8]) );
	inv_0 U89 ( .x(n51), .a(B[6]) );
	aoi21_1 U9 ( .x(n121), .a(A[26]), .b(n69), .c(n122) );
	oa22_3 U91 ( .x(n16), .a(A[13]), .b(n53), .c(A[12]), .d(n52) );
	oa22_1 U92 ( .x(n17), .a(B[9]), .b(n55), .c(B[10]), .d(n54) );
	oa22_1 U93 ( .x(n18), .a(A[6]), .b(n51), .c(A[7]), .d(n49) );
	ao21_3 U94 ( .x(n19), .a(A[20]), .b(n58), .c(n104) );
	inv_2 U95 ( .x(n62), .a(B[15]) );
	nor2i_1 U96 ( .x(n118), .a(A[24]), .b(B[24]) );
	buf_3 U98 ( .x(n20), .a(B[1]) );
	inv_2 U99 ( .x(n24), .a(B[3]) );

endmodule


module EX_DW01_cmp2_32_2 (  A, B, LEQ, TC, LT_LE, GE_GT );

input  LEQ, TC;
input [31:0] A, B;
output  LT_LE, GE_GT;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n15, n16, n17, n18, n19, n20,
	n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
	n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
	n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
	n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
	n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
	n91, n92, n93, n94, n95, n96, n97, n98, n99;


	inv_2 U10 ( .x(n18), .a(A[23]) );
	nand2i_2 U100 ( .x(n48), .a(A[24]), .b(B[24]) );
	inv_0 U101 ( .x(n68), .a(B[17]) );
	nor2i_0 U102 ( .x(n129), .a(B[5]), .b(A[5]) );
	inv_0 U103 ( .x(n95), .a(A[0]) );
	nand2i_0 U104 ( .x(n125), .a(B[3]), .b(A[3]) );
	nand2i_0 U105 ( .x(n34), .a(A[3]), .b(B[3]) );
	nand2i_0 U106 ( .x(n100), .a(B[7]), .b(A[7]) );
	nor2i_0 U107 ( .x(n24), .a(A[8]), .b(B[8]) );
	nand2i_0 U108 ( .x(n39), .a(A[8]), .b(B[8]) );
	inv_0 U109 ( .x(n38), .a(B[9]) );
	inv_2 U11 ( .x(n17), .a(A[25]) );
	oai22_1 U110 ( .x(n76), .a(B[22]), .b(n72), .c(B[21]), .d(n71) );
	nor2i_0 U111 ( .x(n108), .a(B[21]), .b(A[21]) );
	oai22_1 U112 ( .x(n67), .a(B[15]), .b(n42), .c(B[16]), .d(n66) );
	aoi22_1 U113 ( .x(n117), .a(B[16]), .b(n66), .c(B[17]), .d(n93) );
	nand2i_0 U114 ( .x(n118), .a(B[14]), .b(A[14]) );
	aoi22_1 U115 ( .x(n41), .a(B[15]), .b(n42), .c(B[14]), .d(n43) );
	inv_0 U116 ( .x(n90), .a(B[13]) );
	nand2i_0 U117 ( .x(n119), .a(B[13]), .b(A[13]) );
	oai22_1 U118 ( .x(n121), .a(B[11]), .b(n92), .c(B[12]), .d(n91) );
	inv_0 U119 ( .x(n89), .a(B[12]) );
	nand3_2 U12 ( .x(n73), .a(n105), .b(n106), .c(n107) );
	nor2i_0 U120 ( .x(n22), .a(A[6]), .b(B[6]) );
	nand2i_0 U121 ( .x(n140), .a(A[6]), .b(B[6]) );
	aoi22_1 U122 ( .x(n131), .a(B[10]), .b(n97), .c(B[11]), .d(n92) );
	oai22_1 U123 ( .x(n40), .a(B[10]), .b(n97), .c(B[9]), .d(n96) );
	and4i_4 U124 ( .x(n55), .a(n59), .b(n56), .c(n57), .d(n58) );
	nand3i_5 U125 ( .x(n47), .a(n73), .b(n74), .c(n75) );
	nand2i_4 U126 ( .x(n86), .a(n87), .b(n88) );
	nand4i_4 U127 ( .x(n32), .a(n24), .b(n98), .c(n99), .d(n100) );
	oai211_4 U128 ( .x(n87), .a(n41), .b(n67), .c(n117), .d(n16) );
	nand2i_4 U129 ( .x(n59), .a(n132), .b(n133) );
	nand2i_2 U13 ( .x(n106), .a(B[26]), .b(A[26]) );
	nand2_2 U130 ( .x(n132), .a(n15), .b(n131) );
	nand4_1 U131 ( .x(n61), .a(n135), .b(n136), .c(n134), .d(n137) );
	nand2i_4 U132 ( .x(n136), .a(n119), .b(n133) );
	nand2i_4 U133 ( .x(n135), .a(n120), .b(n133) );
	nand2i_6 U134 ( .x(n105), .a(B[27]), .b(A[27]) );
	nand2i_2 U14 ( .x(n107), .a(B[28]), .b(A[28]) );
	nand2i_2 U15 ( .x(n122), .a(B[18]), .b(A[18]) );
	inv_2 U16 ( .x(n91), .a(A[12]) );
	inv_2 U17 ( .x(n92), .a(A[11]) );
	nand3_1 U18 ( .x(n35), .a(n125), .b(n94), .c(B[2]) );
	inv_2 U19 ( .x(n94), .a(A[2]) );
	and4i_1 U20 ( .x(n31), .a(n25), .b(n125), .c(n126), .d(n127) );
	nand2i_2 U21 ( .x(n126), .a(B[2]), .b(A[2]) );
	nand2i_0 U22 ( .x(n127), .a(B[4]), .b(A[4]) );
	nor2i_1 U23 ( .x(n25), .a(n26), .b(n27) );
	inv_2 U24 ( .x(n26), .a(B[0]) );
	nand2i_2 U25 ( .x(n30), .a(n95), .b(n142) );
	nand2i_2 U26 ( .x(n142), .a(A[1]), .b(B[1]) );
	inv_2 U27 ( .x(n27), .a(n142) );
	nand2i_2 U28 ( .x(n29), .a(B[1]), .b(A[1]) );
	inv_2 U29 ( .x(n97), .a(A[10]) );
	inv_2 U30 ( .x(n96), .a(A[9]) );
	nor2i_1 U31 ( .x(n23), .a(A[5]), .b(B[5]) );
	oai211_1 U32 ( .x(n98), .a(n22), .b(n23), .c(n140), .d(n141) );
	inv_2 U33 ( .x(n80), .a(B[19]) );
	inv_2 U34 ( .x(n79), .a(B[18]) );
	inv_2 U35 ( .x(n93), .a(A[17]) );
	inv_2 U36 ( .x(n43), .a(A[14]) );
	nor3i_1 U37 ( .x(n84), .a(n116), .b(n49), .c(n46) );
	nor2_0 U38 ( .x(n49), .a(n47), .b(n50) );
	nor2_0 U39 ( .x(n46), .a(n47), .b(n48) );
	aoi21_1 U40 ( .x(n83), .a(n108), .b(n115), .c(n112) );
	inv_2 U41 ( .x(n115), .a(n54) );
	oai33_1 U42 ( .x(n112), .a(n113), .b(A[27]), .c(n70), .d(n113), .e(n114),
		.f(n103) );
	inv_2 U43 ( .x(n113), .a(n107) );
	inv_2 U44 ( .x(n70), .a(B[27]) );
	nor2i_1 U45 ( .x(n109), .a(B[20]), .b(A[20]) );
	nor2i_1 U46 ( .x(n111), .a(B[23]), .b(A[23]) );
	nor2i_1 U47 ( .x(n110), .a(B[22]), .b(A[22]) );
	inv_0 U48 ( .x(n71), .a(A[21]) );
	inv_0 U49 ( .x(n72), .a(A[22]) );
	nand2i_2 U50 ( .x(n54), .a(n76), .b(n77) );
	nand3_1 U51 ( .x(n124), .a(n16), .b(n68), .c(A[17]) );
	nand2i_2 U52 ( .x(n123), .a(n122), .b(n16) );
	nand3i_1 U53 ( .x(n53), .a(n44), .b(n123), .c(n124) );
	nand2i_2 U54 ( .x(n52), .a(B[20]), .b(A[20]) );
	nand2i_2 U55 ( .x(n137), .a(n118), .b(n133) );
	nor2i_1 U56 ( .x(n102), .a(A[30]), .b(B[30]) );
	inv_2 U57 ( .x(n62), .a(B[30]) );
	inv_2 U58 ( .x(n63), .a(B[31]) );
	oai22_1 U59 ( .x(n64), .a(A[31]), .b(n63), .c(A[30]), .d(n62) );
	nand2i_2 U6 ( .x(n103), .a(A[26]), .b(B[26]) );
	nor2i_1 U60 ( .x(n101), .a(A[29]), .b(B[29]) );
	aoi22_1 U61 ( .x(n134), .a(n101), .b(n85), .c(n102), .d(n85) );
	nand2_2 U62 ( .x(n120), .a(n15), .b(n121) );
	aoi211_1 U63 ( .x(n58), .a(n128), .b(n130), .c(n28), .d(n33) );
	nor2i_1 U64 ( .x(n128), .a(B[4]), .b(A[4]) );
	inv_2 U65 ( .x(n130), .a(n32) );
	inv_2 U66 ( .x(n99), .a(n40) );
	and4i_1 U67 ( .x(n28), .a(n32), .b(n29), .c(n30), .d(n31) );
	aoi211_1 U68 ( .x(n33), .a(n34), .b(n35), .c(n36), .d(n32) );
	inv_2 U69 ( .x(n36), .a(n127) );
	nor2i_2 U7 ( .x(n45), .a(A[25]), .b(B[25]) );
	oaoi211_1 U70 ( .x(n37), .a(A[9]), .b(n38), .c(n39), .d(n40) );
	aoi21_1 U71 ( .x(n57), .a(n129), .b(n130), .c(n37) );
	nand2i_2 U72 ( .x(n56), .a(n19), .b(n130) );
	nor2_1 U73 ( .x(n19), .a(n20), .b(n21) );
	inv_2 U74 ( .x(n20), .a(n140) );
	inv_2 U75 ( .x(n21), .a(n141) );
	inv_4 U76 ( .x(n88), .a(n81) );
	nand2i_2 U77 ( .x(n139), .a(B[31]), .b(A[31]) );
	inv_2 U78 ( .x(n85), .a(n64) );
	nand4_1 U79 ( .x(n81), .a(n82), .b(n83), .c(n84), .d(n85) );
	nor2i_1 U8 ( .x(n104), .a(A[24]), .b(B[24]) );
	nor3i_1 U80 ( .x(n51), .a(n52), .b(n53), .c(n54) );
	inv_2 U81 ( .x(n66), .a(A[16]) );
	inv_0 U82 ( .x(n42), .a(A[15]) );
	nor3i_2 U83 ( .x(LT_LE), .a(n60), .b(n55), .c(n61) );
	inv_5 U84 ( .x(n133), .a(n86) );
	oa22_1 U85 ( .x(n15), .a(A[13]), .b(n90), .c(A[12]), .d(n89) );
	oa22_2 U86 ( .x(n16), .a(A[19]), .b(n80), .c(A[18]), .d(n79) );
	inv_2 U87 ( .x(n69), .a(A[28]) );
	aoi22_1 U88 ( .x(n116), .a(B[28]), .b(n69), .c(n65), .d(B[29]) );
	inv_2 U89 ( .x(n65), .a(A[29]) );
	aoi21_1 U9 ( .x(n75), .a(n104), .b(n50), .c(n45) );
	inv_0 U90 ( .x(n114), .a(n105) );
	nand4i_1 U91 ( .x(n74), .a(n18), .b(n50), .c(n48), .d(n78) );
	inv_5 U92 ( .x(n78), .a(B[23]) );
	inv_7 U93 ( .x(n77), .a(n47) );
	nor2i_1 U94 ( .x(n44), .a(A[19]), .b(B[19]) );
	oai21_1 U95 ( .x(n138), .a(n51), .b(n81), .c(n139) );
	nand2i_0 U96 ( .x(n141), .a(A[7]), .b(B[7]) );
	aoi21_3 U97 ( .x(n60), .a(n133), .b(n67), .c(n138) );
	nand2_5 U98 ( .x(n50), .a(n17), .b(B[25]) );
	aoi222_1 U99 ( .x(n82), .a(n109), .b(n115), .c(n111), .d(n77), .e(n110),
		.f(n77) );

endmodule


module EX_DW01_cmp2_32_4_test_1 (  A, B, LEQ, TC, LT_LE, GE_GT );

input  LEQ, TC;
input [31:0] A, B;
output  LT_LE, GE_GT;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n128, n129, n130, n131, n132, n133, n134, n135, n136,
	n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
	n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
	n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
	n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
	n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
	n71, n72, n73, n74, n75, n76, n77, n79, n80, n81, n82, n83, n84, n85,
	n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	aoi22_1 U10 ( .x(n116), .a(A[25]), .b(n59), .c(n115), .d(n117) );
	inv_2 U101 ( .x(n27), .a(A[20]) );
	inv_2 U102 ( .x(n16), .a(n47) );
	inv_2 U103 ( .x(n47), .a(B[1]) );
	buf_3 U104 ( .x(n17), .a(B[3]) );
	inv_2 U105 ( .x(n18), .a(n84) );
	inv_2 U106 ( .x(n84), .a(A[30]) );
	oai22_1 U107 ( .x(n23), .a(B[17]), .b(n24), .c(B[18]), .d(n25) );
	aoi22_1 U108 ( .x(n97), .a(B[16]), .b(n61), .c(B[17]), .d(n24) );
	oai22_1 U109 ( .x(n120), .a(B[30]), .b(n84), .c(B[29]), .d(n85) );
	inv_2 U11 ( .x(n119), .a(n131) );
	aoi22_1 U110 ( .x(n26), .a(B[20]), .b(n27), .c(B[21]), .d(n28) );
	nor2i_2 U111 ( .x(n21), .a(A[20]), .b(B[20]) );
	oai22_1 U112 ( .x(n141), .a(A[8]), .b(n55), .c(A[9]), .d(n54) );
	nor2i_0 U113 ( .x(n29), .a(A[8]), .b(B[8]) );
	ao222_3 U114 ( .x(n19), .a(A[0]), .b(n147), .c(n147), .d(n44), .e(n94),
		.f(n147) );
	oai22_1 U115 ( .x(n135), .a(B[11]), .b(n87), .c(B[12]), .d(n86) );
	nand2i_0 U116 ( .x(n76), .a(A[11]), .b(B[11]) );
	nand2i_0 U117 ( .x(n91), .a(A[3]), .b(n17) );
	inv_0 U118 ( .x(n40), .a(A[3]) );
	inv_0 U119 ( .x(n49), .a(B[0]) );
	aoi21_1 U12 ( .x(n118), .a(A[26]), .b(n64), .c(n119) );
	oai22_1 U120 ( .x(n77), .a(A[6]), .b(n43), .c(A[7]), .d(n42) );
	aoi211_1 U121 ( .x(n37), .a(A[7]), .b(n42), .c(n29), .d(n56) );
	nand2i_2 U122 ( .x(n32), .a(A[18]), .b(B[18]) );
	oai22_1 U123 ( .x(n56), .a(B[10]), .b(n53), .c(B[9]), .d(n52) );
	inv_0 U124 ( .x(n54), .a(B[9]) );
	aoi21_1 U125 ( .x(n111), .a(A[13]), .b(n50), .c(n23) );
	nor2_5 U126 ( .x(LT_LE), .a(n19), .b(n20) );
	aoi21_6 U127 ( .x(n31), .a(n32), .b(n33), .c(n34) );
	nor2i_5 U128 ( .x(n98), .a(n99), .b(n34) );
	nand2i_4 U129 ( .x(n101), .a(A[27]), .b(B[27]) );
	nor3i_5 U130 ( .x(n74), .a(n106), .b(n67), .c(n31) );
	nand2i_4 U131 ( .x(n110), .a(n92), .b(n140) );
	nand3i_5 U132 ( .x(n20), .a(n35), .b(n128), .c(n129) );
	nand2i_6 U134 ( .x(n82), .a(B[2]), .b(A[2]) );
	nand2_4 U135 ( .x(n72), .a(n98), .b(n145) );
	nand3i_5 U136 ( .x(n108), .a(n107), .b(n109), .c(n110) );
	nand3i_5 U137 ( .x(n67), .a(n68), .b(n69), .c(n70) );
	nand2i_6 U138 ( .x(n131), .a(B[27]), .b(A[27]) );
	inv_0 U139 ( .x(n66), .a(B[29]) );
	inv_2 U14 ( .x(n144), .a(n132) );
	and4_5 U140 ( .x(n147), .a(n148), .b(n79), .c(n80), .d(n81) );
	inv_3 U141 ( .x(n148), .a(n39) );
	nand4i_2 U142 ( .x(n39), .a(n71), .b(n72), .c(n73), .d(n74) );
	nor2_2 U143 ( .x(n80), .a(n38), .b(n77) );
	nand2i_0 U144 ( .x(n132), .a(B[28]), .b(A[28]) );
	inv_0 U145 ( .x(n65), .a(B[28]) );
	nor2i_0 U146 ( .x(n100), .a(B[26]), .b(A[26]) );
	nand2i_4 U147 ( .x(n134), .a(A[24]), .b(B[24]) );
	nand4i_1 U15 ( .x(n123), .a(n144), .b(n118), .c(n116), .d(n133) );
	nand2i_2 U16 ( .x(n113), .a(B[14]), .b(A[14]) );
	inv_2 U17 ( .x(n86), .a(A[12]) );
	inv_2 U18 ( .x(n87), .a(A[11]) );
	nand2i_0 U19 ( .x(n92), .a(A[2]), .b(B[2]) );
	nand2i_2 U20 ( .x(n109), .a(n91), .b(n140) );
	inv_2 U21 ( .x(n140), .a(n44) );
	inv_2 U22 ( .x(n41), .a(A[4]) );
	inv_2 U23 ( .x(n45), .a(B[4]) );
	oai22_1 U24 ( .x(n107), .a(A[4]), .b(n45), .c(A[5]), .d(n46) );
	inv_0 U25 ( .x(n51), .a(B[12]) );
	nand2_2 U26 ( .x(n75), .a(n137), .b(n141) );
	nor2i_0 U27 ( .x(n30), .a(B[10]), .b(A[10]) );
	nand2i_2 U28 ( .x(n33), .a(A[19]), .b(B[19]) );
	nand3_1 U29 ( .x(n70), .a(n131), .b(n100), .c(n132) );
	nand2i_2 U30 ( .x(n69), .a(n101), .b(n132) );
	oai22_1 U32 ( .x(n68), .a(A[29]), .b(n66), .c(A[28]), .d(n65) );
	nand2i_2 U33 ( .x(n130), .a(B[31]), .b(A[31]) );
	nor2i_1 U34 ( .x(n96), .a(B[30]), .b(n18) );
	inv_0 U35 ( .x(n114), .a(n63) );
	inv_2 U36 ( .x(n61), .a(A[16]) );
	inv_5 U37 ( .x(n62), .a(A[15]) );
	oai22_1 U38 ( .x(n63), .a(B[15]), .b(n62), .c(B[16]), .d(n61) );
	nand2i_2 U39 ( .x(n142), .a(A[14]), .b(B[14]) );
	aoai211_1 U40 ( .x(n145), .a(n143), .b(n142), .c(n63), .d(n97) );
	or3i_2 U41 ( .x(n34), .a(n60), .b(n21), .c(n22) );
	inv_2 U42 ( .x(n25), .a(A[18]) );
	inv_2 U43 ( .x(n24), .a(A[17]) );
	inv_2 U44 ( .x(n99), .a(n23) );
	inv_2 U45 ( .x(n105), .a(n134) );
	nand2i_2 U46 ( .x(n117), .a(A[25]), .b(B[25]) );
	inv_2 U47 ( .x(n104), .a(n117) );
	nor2_1 U48 ( .x(n103), .a(n104), .b(n105) );
	inv_2 U49 ( .x(n88), .a(A[23]) );
	aoi22_1 U50 ( .x(n102), .a(B[23]), .b(n88), .c(B[22]), .d(n57) );
	oai22_1 U51 ( .x(n58), .a(B[21]), .b(n28), .c(B[22]), .d(n57) );
	inv_0 U52 ( .x(n28), .a(A[21]) );
	inv_2 U53 ( .x(n57), .a(A[22]) );
	inv_2 U54 ( .x(n60), .a(n58) );
	inv_0 U55 ( .x(n64), .a(B[26]) );
	inv_2 U56 ( .x(n124), .a(n130) );
	inv_2 U57 ( .x(n122), .a(n67) );
	aoi211_1 U58 ( .x(n121), .a(n122), .b(n123), .c(n124), .d(n120) );
	and4i_1 U59 ( .x(n112), .a(n34), .b(n113), .c(n114), .d(n111) );
	nand2_2 U60 ( .x(n136), .a(n15), .b(n135) );
	aoai211_1 U61 ( .x(n146), .a(n136), .b(n112), .c(n39), .d(n121) );
	nand2i_2 U62 ( .x(n106), .a(A[31]), .b(B[31]) );
	inv_2 U63 ( .x(n126), .a(n106) );
	nand2i_2 U64 ( .x(n125), .a(n126), .b(n73) );
	inv_0 U65 ( .x(n53), .a(A[10]) );
	inv_0 U66 ( .x(n52), .a(A[9]) );
	inv_2 U67 ( .x(n137), .a(n56) );
	inv_0 U68 ( .x(n89), .a(A[5]) );
	inv_0 U69 ( .x(n90), .a(A[6]) );
	nor2i_1 U7 ( .x(n22), .a(A[19]), .b(B[19]) );
	oai22_1 U70 ( .x(n139), .a(B[6]), .b(n90), .c(B[5]), .d(n89) );
	nand2_2 U71 ( .x(n36), .a(n138), .b(n139) );
	aoi21_2 U72 ( .x(n81), .a(n95), .b(n93), .c(n108) );
	nor2_1 U73 ( .x(n95), .a(n44), .b(n47) );
	nor2i_1 U74 ( .x(n93), .a(n48), .b(n94) );
	inv_2 U75 ( .x(n48), .a(A[1]) );
	inv_2 U76 ( .x(n138), .a(n77) );
	nand4i_1 U77 ( .x(n38), .a(n30), .b(n75), .c(n15), .d(n76) );
	nand2i_2 U79 ( .x(n83), .a(n16), .b(A[1]) );
	inv_2 U8 ( .x(n85), .a(A[29]) );
	nand4i_1 U80 ( .x(n79), .a(n49), .b(n140), .c(n83), .d(n82) );
	oai211_1 U82 ( .x(n71), .a(n26), .b(n58), .c(n102), .d(n103) );
	nand2_2 U83 ( .x(n73), .a(n96), .b(n130) );
	nand2i_2 U84 ( .x(n129), .a(n83), .b(n147) );
	nand2i_2 U85 ( .x(n128), .a(n125), .b(n146) );
	aoi211_1 U86 ( .x(n35), .a(n36), .b(n37), .c(n38), .d(n39) );
	inv_2 U87 ( .x(n94), .a(n82) );
	oai22_1 U88 ( .x(n44), .a(B[4]), .b(n41), .c(n17), .d(n40) );
	nand4i_1 U9 ( .x(n133), .a(B[23]), .b(n117), .c(A[23]), .d(n134) );
	inv_0 U90 ( .x(n50), .a(B[13]) );
	inv_0 U91 ( .x(n46), .a(B[5]) );
	inv_2 U92 ( .x(n59), .a(B[25]) );
	inv_2 U93 ( .x(n42), .a(B[7]) );
	inv_0 U94 ( .x(n55), .a(B[8]) );
	inv_0 U95 ( .x(n43), .a(B[6]) );
	oa22_2 U97 ( .x(n15), .a(A[12]), .b(n51), .c(A[13]), .d(n50) );
	nand2i_2 U98 ( .x(n143), .a(A[15]), .b(B[15]) );
	nor2i_1 U99 ( .x(n115), .a(A[24]), .b(B[24]) );

endmodule


module EX_DW01_cmp2_32_1 (  A, B, LEQ, TC, LT_LE, GE_GT );

input  LEQ, TC;
input [31:0] A, B;
output  LT_LE, GE_GT;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n15, n16, n17, n18, n19, n20, n21, n22,
	n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
	n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
	n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
	n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
	n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
	n93, n94, n95, n96, n97, n98, n99;


	and4_3 U10 ( .x(n18), .a(A[23]), .b(n85), .c(n84), .d(n81) );
	nand2i_0 U100 ( .x(n103), .a(B[5]), .b(A[5]) );
	nand2i_0 U101 ( .x(n109), .a(A[5]), .b(B[5]) );
	oai22_1 U102 ( .x(n112), .a(A[9]), .b(n87), .c(A[8]), .d(n86) );
	inv_0 U103 ( .x(n88), .a(A[0]) );
	inv_0 U104 ( .x(n32), .a(A[3]) );
	nand2i_0 U105 ( .x(n106), .a(B[3]), .b(A[3]) );
	aoi22_1 U106 ( .x(n102), .a(A[7]), .b(n66), .c(A[8]), .d(n86) );
	oai22_1 U107 ( .x(n67), .a(A[7]), .b(n66), .c(A[6]), .d(n65) );
	inv_0 U108 ( .x(n86), .a(B[8]) );
	inv_0 U109 ( .x(n87), .a(B[9]) );
	inv_2 U11 ( .x(n81), .a(B[23]) );
	oai22_1 U110 ( .x(n60), .a(B[21]), .b(n57), .c(B[22]), .d(n56) );
	nand2i_0 U111 ( .x(n97), .a(A[21]), .b(B[21]) );
	inv_0 U112 ( .x(n27), .a(B[16]) );
	nor2i_0 U113 ( .x(n37), .a(B[16]), .b(A[16]) );
	inv_0 U114 ( .x(n35), .a(B[14]) );
	aoi22_1 U115 ( .x(n98), .a(A[13]), .b(n71), .c(A[14]), .d(n35) );
	oai22_1 U116 ( .x(n72), .a(A[13]), .b(n71), .c(A[12]), .d(n25) );
	nand2i_0 U117 ( .x(n104), .a(B[6]), .b(A[6]) );
	inv_0 U118 ( .x(n65), .a(B[6]) );
	aoi221_1 U119 ( .x(n43), .a(n111), .b(n112), .c(B[10]), .d(n64), .e(n33) );
	nand3_1 U12 ( .x(n58), .a(n93), .b(n94), .c(n95) );
	oai22_1 U120 ( .x(n78), .a(B[10]), .b(n64), .c(B[9]), .d(n63) );
	nor3i_5 U121 ( .x(n45), .a(n46), .b(n47), .c(n48) );
	aoi21_3 U122 ( .x(LT_LE), .a(n49), .b(n50), .c(n51) );
	or3i_5 U123 ( .x(n48), .a(n80), .b(n78), .c(n79) );
	or3i_4 U124 ( .x(n125), .a(n135), .b(n30), .c(n105) );
	nand2i_4 U125 ( .x(n128), .a(n108), .b(n135) );
	nand2i_4 U126 ( .x(n127), .a(n109), .b(n135) );
	inv_7 U127 ( .x(n135), .a(n48) );
	nand2i_5 U128 ( .x(n124), .a(n121), .b(n125) );
	nand2i_5 U129 ( .x(n76), .a(n26), .b(n114) );
	nand2i_2 U13 ( .x(n94), .a(B[26]), .b(A[26]) );
	inv_6 U130 ( .x(n114), .a(n70) );
	nand2i_5 U131 ( .x(n59), .a(n60), .b(n17) );
	inv_10 U132 ( .x(n57), .a(A[21]) );
	nand2i_2 U14 ( .x(n95), .a(B[28]), .b(A[28]) );
	nor2i_0 U15 ( .x(n33), .a(B[11]), .b(A[11]) );
	inv_0 U16 ( .x(n71), .a(B[13]) );
	nand2i_0 U17 ( .x(n139), .a(B[11]), .b(A[11]) );
	aoai211_1 U18 ( .x(n140), .a(n139), .b(n15), .c(n72), .d(n98) );
	oai22_1 U19 ( .x(n34), .a(A[14]), .b(n35), .c(A[15]), .d(n28) );
	inv_2 U20 ( .x(n24), .a(A[18]) );
	nor2i_1 U21 ( .x(n36), .a(B[17]), .b(A[17]) );
	or3i_2 U22 ( .x(n70), .a(n22), .b(n36), .c(n37) );
	inv_2 U23 ( .x(n28), .a(B[15]) );
	aoi22_1 U24 ( .x(n26), .a(A[16]), .b(n27), .c(A[15]), .d(n28) );
	inv_0 U25 ( .x(n56), .a(A[22]) );
	aoi22_1 U26 ( .x(n22), .a(n24), .b(B[18]), .c(n23), .d(B[19]) );
	inv_2 U27 ( .x(n23), .a(A[19]) );
	inv_2 U28 ( .x(n19), .a(A[20]) );
	inv_2 U29 ( .x(n61), .a(B[20]) );
	inv_0 U30 ( .x(n68), .a(B[19]) );
	nand2i_0 U31 ( .x(n101), .a(B[17]), .b(A[17]) );
	nand2i_2 U32 ( .x(n100), .a(B[18]), .b(A[18]) );
	nand2i_2 U33 ( .x(n89), .a(B[29]), .b(A[29]) );
	nand2_2 U34 ( .x(n105), .a(n106), .b(n107) );
	inv_2 U35 ( .x(n31), .a(A[2]) );
	aoi22_1 U36 ( .x(n30), .a(B[2]), .b(n31), .c(B[3]), .d(n32) );
	nand3i_1 U37 ( .x(n121), .a(n118), .b(n122), .c(n123) );
	inv_2 U38 ( .x(n119), .a(n95) );
	inv_2 U39 ( .x(n55), .a(B[27]) );
	nand2i_0 U40 ( .x(n122), .a(n96), .b(n75) );
	nand2i_0 U41 ( .x(n123), .a(n97), .b(n75) );
	nor2_1 U42 ( .x(n38), .a(n39), .b(n40) );
	nor3_2 U43 ( .x(n17), .a(n58), .b(n18), .c(n16) );
	nand2i_2 U44 ( .x(n40), .a(A[22]), .b(B[22]) );
	nor2i_1 U45 ( .x(n110), .a(B[23]), .b(A[23]) );
	nand2i_2 U46 ( .x(n108), .a(A[4]), .b(B[4]) );
	aoi21_1 U47 ( .x(n130), .a(n131), .b(n17), .c(n129) );
	inv_2 U48 ( .x(n131), .a(n84) );
	nand2i_2 U49 ( .x(n84), .a(A[24]), .b(B[24]) );
	oai22_1 U50 ( .x(n129), .a(A[29]), .b(n83), .c(A[28]), .d(n82) );
	inv_2 U51 ( .x(n83), .a(B[29]) );
	inv_2 U52 ( .x(n82), .a(B[28]) );
	nand2i_2 U53 ( .x(n85), .a(A[25]), .b(B[25]) );
	inv_2 U54 ( .x(n134), .a(n85) );
	aoi21_1 U55 ( .x(n133), .a(n134), .b(n17), .c(n54) );
	nand3i_2 U56 ( .x(n77), .a(n34), .b(n114), .c(n140) );
	nor2i_1 U57 ( .x(n42), .a(n43), .b(n44) );
	nand3i_0 U58 ( .x(n44), .a(n72), .b(n113), .c(n114) );
	inv_2 U59 ( .x(n113), .a(n34) );
	nand2i_2 U6 ( .x(n96), .a(n20), .b(B[20]) );
	oai31_2 U60 ( .x(n47), .a(n88), .b(B[0]), .c(n29), .d(n117) );
	nor2i_1 U61 ( .x(n29), .a(B[1]), .b(A[1]) );
	nand2i_2 U62 ( .x(n117), .a(B[1]), .b(A[1]) );
	aoi211_1 U63 ( .x(n46), .a(A[2]), .b(n62), .c(n115), .d(n116) );
	inv_2 U64 ( .x(n62), .a(B[2]) );
	inv_2 U65 ( .x(n115), .a(n107) );
	nand2i_2 U66 ( .x(n107), .a(B[4]), .b(A[4]) );
	inv_2 U67 ( .x(n116), .a(n106) );
	nand4i_1 U68 ( .x(n73), .a(n74), .b(n75), .c(n76), .d(n77) );
	aoai211_1 U69 ( .x(n74), .a(n100), .b(n101), .c(n69), .d(n99) );
	nand2i_2 U7 ( .x(n91), .a(A[26]), .b(B[26]) );
	inv_5 U70 ( .x(n75), .a(n59) );
	inv_2 U71 ( .x(n80), .a(n73) );
	aoai211_1 U72 ( .x(n79), .a(n103), .b(n104), .c(n67), .d(n102) );
	inv_0 U73 ( .x(n64), .a(A[10]) );
	inv_0 U74 ( .x(n63), .a(A[9]) );
	inv_2 U75 ( .x(n111), .a(n78) );
	nand2i_2 U76 ( .x(n137), .a(B[31]), .b(A[31]) );
	inv_2 U77 ( .x(n138), .a(n54) );
	nand2i_2 U78 ( .x(n136), .a(n89), .b(n138) );
	nand2i_2 U79 ( .x(n90), .a(B[30]), .b(A[30]) );
	nor2i_0 U8 ( .x(n41), .a(A[25]), .b(B[25]) );
	inv_2 U80 ( .x(n52), .a(B[30]) );
	inv_2 U81 ( .x(n53), .a(B[31]) );
	oai22_1 U82 ( .x(n54), .a(A[31]), .b(n53), .c(A[30]), .d(n52) );
	oai211_1 U83 ( .x(n51), .a(n54), .b(n90), .c(n136), .d(n137) );
	and4i_3 U84 ( .x(n50), .a(n124), .b(n127), .c(n128), .d(n126) );
	aoi21_1 U85 ( .x(n126), .a(n110), .b(n17), .c(n38) );
	aoi211_1 U86 ( .x(n49), .a(n135), .b(n67), .c(n45), .d(n132) );
	inv_0 U87 ( .x(n66), .a(B[7]) );
	oai211_1 U88 ( .x(n132), .a(n42), .b(n21), .c(n133), .d(n130) );
	nand2_2 U89 ( .x(n15), .a(n25), .b(A[12]) );
	nor2i_1 U9 ( .x(n92), .a(A[24]), .b(B[24]) );
	ao21_3 U90 ( .x(n16), .a(n92), .b(n85), .c(n41) );
	inv_0 U91 ( .x(n39), .a(n17) );
	oai33_1 U92 ( .x(n118), .a(n119), .b(A[27]), .c(n55), .d(n119), .e(n120),
		.f(n91) );
	inv_0 U93 ( .x(n120), .a(n93) );
	nand2i_4 U94 ( .x(n93), .a(B[27]), .b(A[27]) );
	inv_2 U95 ( .x(n20), .a(n19) );
	nand4i_1 U96 ( .x(n21), .a(n74), .b(n75), .c(n76), .d(n77) );
	aoi22_1 U97 ( .x(n99), .a(n20), .b(n61), .c(A[19]), .d(n68) );
	inv_2 U98 ( .x(n69), .a(n22) );
	inv_0 U99 ( .x(n25), .a(B[12]) );

endmodule


module EX_DW01_sub_32_2_test_1 (  A, B, CI, DIFF, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] DIFF;

wire n100, n101, n102, n103, n104, n105, n108, n109, n110, n111, n112, n113,
	n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
	n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
	n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
	n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
	n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
	n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185,
	n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
	n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
	n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
	n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
	n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
	n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
	n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
	n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
	n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
	n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
	n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
	n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
	n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
	n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
	n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
	n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
	n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
	n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
	n92, n93, n94, n95, n96, n97, n98, n99;


	inv_2 U10 ( .x(n191), .a(n59) );
	inv_2 U100 ( .x(n218), .a(n318) );
	oai21_1 U101 ( .x(n214), .a(n121), .b(n51), .c(n250) );
	inv_0 U102 ( .x(n171), .a(n284) );
	nor2_1 U103 ( .x(n169), .a(n170), .b(n171) );
	nand2i_2 U104 ( .x(n333), .a(B[14]), .b(A[14]) );
	inv_2 U105 ( .x(n173), .a(n333) );
	oai21_1 U106 ( .x(n228), .a(n82), .b(n50), .c(n141) );
	nor2_1 U107 ( .x(n167), .a(n168), .b(n311) );
	inv_2 U108 ( .x(n168), .a(n200) );
	inv_2 U109 ( .x(n311), .a(n330) );
	nor2_1 U110 ( .x(n79), .a(A[16]), .b(n80) );
	inv_2 U111 ( .x(n360), .a(n329) );
	aoi211_1 U112 ( .x(n190), .a(n191), .b(n192), .c(n193), .d(n194) );
	oai211_2 U113 ( .x(n331), .a(n190), .b(n255), .c(n332), .d(n328) );
	nand2i_2 U114 ( .x(n147), .a(B[21]), .b(A[21]) );
	inv_2 U115 ( .x(n337), .a(n147) );
	nand2i_2 U116 ( .x(n300), .a(B[21]), .b(n299) );
	inv_2 U117 ( .x(n257), .a(A[21]) );
	nand2i_2 U118 ( .x(n298), .a(n257), .b(n299) );
	nor2i_0 U119 ( .x(n148), .a(A[22]), .b(B[22]) );
	inv_5 U12 ( .x(n175), .a(n247) );
	nand2i_2 U120 ( .x(n342), .a(B[25]), .b(A[25]) );
	inv_2 U121 ( .x(n304), .a(n342) );
	inv_2 U122 ( .x(n302), .a(n240) );
	nand2i_2 U123 ( .x(n303), .a(A[25]), .b(B[25]) );
	exor2_1 U124 ( .x(DIFF[3]), .a(n221), .b(n153) );
	oai21_1 U125 ( .x(n221), .a(n161), .b(n352), .c(n315) );
	inv_2 U126 ( .x(n154), .a(B[3]) );
	exor2_1 U127 ( .x(DIFF[2]), .a(n226), .b(n159) );
	aoai211_1 U128 ( .x(n226), .a(B[1]), .b(n186), .c(n276), .d(n232) );
	nor2_1 U129 ( .x(n159), .a(n160), .b(n161) );
	inv_2 U13 ( .x(n246), .a(n81) );
	inv_2 U130 ( .x(n160), .a(n315) );
	inv_2 U131 ( .x(n161), .a(n277) );
	inv_2 U132 ( .x(n352), .a(n226) );
	exor2_1 U133 ( .x(DIFF[6]), .a(n216), .b(n125) );
	exor2_1 U134 ( .x(DIFF[12]), .a(n229), .b(n177) );
	nor2_1 U135 ( .x(n156), .a(n157), .b(n158) );
	exor2_1 U136 ( .x(DIFF[27]), .a(n223), .b(n156) );
	exor2_1 U137 ( .x(DIFF[11]), .a(n230), .b(n180) );
	exnor2_1 U138 ( .x(DIFF[20]), .a(n209), .b(n272) );
	exor2_1 U139 ( .x(DIFF[14]), .a(n228), .b(n172) );
	nor2i_1 U14 ( .x(n283), .a(n284), .b(n173) );
	exnor2_1 U140 ( .x(DIFF[13]), .a(n50), .b(n174) );
	exor2_1 U141 ( .x(DIFF[10]), .a(n231), .b(n183) );
	exnor2_1 U142 ( .x(DIFF[22]), .a(n146), .b(n270) );
	nor3i_1 U143 ( .x(n146), .a(n147), .b(n144), .c(n112) );
	exnor2_1 U144 ( .x(n270), .a(A[22]), .b(B[22]) );
	exor2_1 U145 ( .x(DIFF[5]), .a(n217), .b(n128) );
	exnor2_1 U146 ( .x(DIFF[19]), .a(n162), .b(n203) );
	nor2_0 U147 ( .x(n162), .a(n88), .b(n163) );
	inv_2 U148 ( .x(n163), .a(n328) );
	exnor2_1 U149 ( .x(DIFF[4]), .a(n218), .b(n131) );
	oai21_1 U15 ( .x(n285), .a(n246), .b(n249), .c(n283) );
	inv_2 U150 ( .x(n198), .a(n310) );
	exnor2_1 U151 ( .x(DIFF[18]), .a(n195), .b(n273) );
	inv_2 U152 ( .x(n347), .a(n309) );
	inv_2 U153 ( .x(n157), .a(n344) );
	exnor2_1 U154 ( .x(DIFF[8]), .a(n51), .b(n120) );
	inv_2 U155 ( .x(n121), .a(n245) );
	mux2i_1 U156 ( .x(DIFF[1]), .d0(n185), .sl(n276), .d1(n275) );
	exor2_1 U157 ( .x(DIFF[9]), .a(n214), .b(n117) );
	mux2i_1 U158 ( .x(DIFF[17]), .d0(n164), .sl(n199), .d1(n274) );
	inv_4 U159 ( .x(n210), .a(n253) );
	nor2_1 U16 ( .x(n139), .a(n140), .b(n141) );
	exnor2_1 U160 ( .x(n271), .a(A[21]), .b(B[21]) );
	exnor2_1 U161 ( .x(n269), .a(A[23]), .b(B[23]) );
	nand2_2 U162 ( .x(n225), .a(n303), .b(n342) );
	inv_2 U163 ( .x(n239), .a(A[24]) );
	exnor2_1 U164 ( .x(DIFF[25]), .a(n224), .b(n225) );
	exnor2_1 U165 ( .x(n265), .a(B[26]), .b(A[26]) );
	exnor2_1 U166 ( .x(DIFF[21]), .a(n113), .b(n271) );
	inv_2 U168 ( .x(n237), .a(B[28]) );
	inv_2 U169 ( .x(n155), .a(n115) );
	inv_0 U17 ( .x(n280), .a(n233) );
	oa21_2 U170 ( .x(n51), .a(n218), .b(n279), .c(n281) );
	inv_2 U171 ( .x(n248), .a(n84) );
	nand2i_3 U172 ( .x(n325), .a(B[9]), .b(A[9]) );
	inv_5 U173 ( .x(n118), .a(n325) );
	exnor2_3 U175 ( .x(DIFF[28]), .a(n53), .b(n52) );
	inv_2 U176 ( .x(n52), .a(n263) );
	ao21_3 U177 ( .x(n53), .a(n212), .b(n213), .c(n157) );
	nand2i_2 U179 ( .x(n284), .a(B[15]), .b(A[15]) );
	and4_3 U18 ( .x(n57), .a(n277), .b(n110), .c(n278), .d(n115) );
	exnor2_1 U180 ( .x(n267), .a(A[24]), .b(B[24]) );
	nand2i_2 U181 ( .x(n359), .a(B[24]), .b(n303) );
	nand2i_2 U182 ( .x(n240), .a(B[24]), .b(A[24]) );
	exnor2_1 U183 ( .x(n263), .a(A[28]), .b(B[28]) );
	nand2i_2 U184 ( .x(n346), .a(A[28]), .b(n344) );
	nand2i_0 U185 ( .x(n355), .a(A[28]), .b(B[28]) );
	inv_2 U186 ( .x(n54), .a(n250) );
	nor2i_3 U187 ( .x(n98), .a(n100), .b(n99) );
	inv_2 U188 ( .x(n202), .a(n88) );
	nor2_4 U189 ( .x(n254), .a(n166), .b(n88) );
	inv_5 U19 ( .x(n65), .a(n179) );
	nor2i_1 U190 ( .x(n142), .a(n143), .b(n88) );
	nor2i_3 U191 ( .x(n88), .a(n90), .b(n89) );
	nor2i_3 U192 ( .x(n290), .a(n291), .b(n233) );
	inv_0 U193 ( .x(n82), .a(n247) );
	inv_0 U194 ( .x(n55), .a(n313) );
	inv_2 U195 ( .x(n56), .a(n55) );
	nand3_2 U197 ( .x(n296), .a(n57), .b(n63), .c(n290) );
	or3i_2 U20 ( .x(n288), .a(n316), .b(n160), .c(A[3]) );
	nor2_3 U200 ( .x(n259), .a(n58), .b(n118) );
	nor3i_5 U202 ( .x(n63), .a(n81), .b(n64), .c(n241) );
	or3i_2 U203 ( .x(n289), .a(n63), .b(n233), .c(n155) );
	exor2_1 U204 ( .x(n275), .a(B[1]), .b(A[1]) );
	inv_0 U205 ( .x(n186), .a(A[1]) );
	nand2i_2 U207 ( .x(n278), .a(A[1]), .b(B[1]) );
	aoi21_1 U208 ( .x(n153), .a(A[3]), .b(n154), .c(n155) );
	nand2_8 U209 ( .x(n59), .a(A[16]), .b(n80) );
	exnor2_5 U210 ( .x(DIFF[31]), .a(n219), .b(n105) );
	exnor2_1 U211 ( .x(DIFF[24]), .a(n266), .b(n267) );
	aoai211_3 U212 ( .x(n101), .a(n359), .b(n358), .c(n266), .d(n301) );
	aoai211_4 U213 ( .x(n102), .a(n359), .b(n358), .c(n266), .d(n301) );
	aoi21_2 U214 ( .x(n201), .a(A[20]), .b(n202), .c(n142) );
	oai21_2 U215 ( .x(n295), .a(n286), .b(n289), .c(n296) );
	or3i_3 U216 ( .x(n336), .a(n258), .b(n179), .c(n246) );
	nand2_2 U217 ( .x(n261), .a(n242), .b(n243) );
	inv_3 U218 ( .x(n138), .a(n63) );
	inv_0 U219 ( .x(n60), .a(n241) );
	or3i_3 U22 ( .x(n287), .a(n316), .b(n160), .c(n154) );
	inv_2 U220 ( .x(n61), .a(n60) );
	nand2i_2 U221 ( .x(n321), .a(B[4]), .b(A[4]) );
	nand2i_2 U222 ( .x(n291), .a(A[4]), .b(B[4]) );
	nand4_4 U223 ( .x(n241), .a(n242), .b(n243), .c(n244), .d(n245) );
	inv_10 U224 ( .x(n242), .a(n66) );
	buf_2 U225 ( .x(n62), .a(n234) );
	nand2i_2 U226 ( .x(n181), .a(B[11]), .b(A[11]) );
	inv_0 U227 ( .x(n208), .a(n331) );
	aoi21_3 U229 ( .x(n292), .a(n293), .b(n294), .c(n135) );
	ao211_5 U231 ( .x(n357), .a(n197), .b(n97), .c(n95), .d(n96) );
	inv_3 U232 ( .x(n97), .a(n297) );
	nor2i_1 U233 ( .x(n92), .a(A[5]), .b(B[5]) );
	oai21_1 U234 ( .x(n256), .a(A[17]), .b(n165), .c(n194) );
	aoai211_1 U235 ( .x(n310), .a(A[17]), .b(n165), .c(n311), .d(n312) );
	aoi21_1 U236 ( .x(n164), .a(A[17]), .b(n165), .c(n166) );
	nand2_6 U237 ( .x(n64), .a(n294), .b(n65) );
	inv_7 U238 ( .x(n179), .a(n334) );
	nor2_8 U239 ( .x(n66), .a(A[10]), .b(n67) );
	nand2i_2 U24 ( .x(n115), .a(A[3]), .b(B[3]) );
	exnor2_3 U240 ( .x(DIFF[30]), .a(n262), .b(n68) );
	exnor2_1 U241 ( .x(n68), .a(A[30]), .b(n69) );
	inv_0 U242 ( .x(n69), .a(B[30]) );
	nand2i_2 U244 ( .x(n308), .a(A[30]), .b(n309) );
	buf_1 U245 ( .x(n70), .a(n212) );
	inv_2 U246 ( .x(n165), .a(B[17]) );
	exor2_1 U247 ( .x(n274), .a(A[17]), .b(B[17]) );
	nand2i_0 U248 ( .x(n312), .a(A[17]), .b(B[17]) );
	nand2i_2 U249 ( .x(n329), .a(B[17]), .b(A[17]) );
	nand2i_2 U25 ( .x(n277), .a(A[2]), .b(B[2]) );
	nand2i_2 U250 ( .x(n192), .a(A[17]), .b(B[17]) );
	nor2i_2 U251 ( .x(n193), .a(A[17]), .b(B[17]) );
	nand2i_2 U252 ( .x(n314), .a(A[17]), .b(B[17]) );
	exnor2_3 U253 ( .x(DIFF[29]), .a(n75), .b(n71) );
	inv_2 U254 ( .x(n71), .a(n222) );
	exnor2_1 U255 ( .x(n72), .a(n74), .b(n73) );
	inv_2 U256 ( .x(n222), .a(n72) );
	inv_0 U257 ( .x(n73), .a(B[29]) );
	inv_2 U258 ( .x(n74), .a(A[29]) );
	aoai211_1 U259 ( .x(n75), .a(n70), .b(n76), .c(n77), .d(n355) );
	nand2i_3 U26 ( .x(n315), .a(B[2]), .b(A[2]) );
	inv_2 U260 ( .x(n76), .a(n158) );
	and2_1 U261 ( .x(n77), .a(n346), .b(n345) );
	inv_2 U262 ( .x(n211), .a(n355) );
	inv_2 U263 ( .x(n158), .a(n213) );
	inv_2 U265 ( .x(n264), .a(n102) );
	nand2i_2 U266 ( .x(n309), .a(B[29]), .b(A[29]) );
	exnor2_1 U268 ( .x(n272), .a(A[20]), .b(B[20]) );
	nor2i_0 U269 ( .x(n134), .a(B[20]), .b(A[20]) );
	nor2_1 U27 ( .x(n125), .a(n126), .b(n127) );
	inv_0 U270 ( .x(n143), .a(B[20]) );
	nor2i_2 U271 ( .x(n78), .a(n252), .b(n79) );
	inv_0 U272 ( .x(n251), .a(n78) );
	inv_0 U273 ( .x(n200), .a(n79) );
	inv_2 U274 ( .x(n80), .a(B[16]) );
	nor2_8 U275 ( .x(n81), .a(n84), .b(n175) );
	nor2_8 U276 ( .x(n84), .a(A[14]), .b(n85) );
	inv_0 U277 ( .x(n170), .a(n294) );
	aoai211_1 U278 ( .x(n224), .a(B[24]), .b(n239), .c(n266), .d(n240) );
	nand2i_0 U279 ( .x(n86), .a(n295), .b(n292) );
	nand3i_3 U282 ( .x(n219), .a(n189), .b(n351), .c(n350) );
	inv_0 U283 ( .x(n87), .a(B[30]) );
	ao211_5 U284 ( .x(n93), .a(n197), .b(n97), .c(n96), .d(n95) );
	inv_2 U285 ( .x(n90), .a(A[19]) );
	aoai211_3 U286 ( .x(n258), .a(n259), .b(n260), .c(n261), .d(n181) );
	inv_0 U287 ( .x(n184), .a(n242) );
	inv_2 U288 ( .x(n91), .a(n129) );
	inv_0 U289 ( .x(n129), .a(n322) );
	oai21_1 U29 ( .x(n216), .a(n130), .b(n326), .c(n91) );
	inv_2 U290 ( .x(n322), .a(n92) );
	nand2i_4 U291 ( .x(n299), .a(A[22]), .b(B[22]) );
	inv_8 U292 ( .x(n255), .a(A[18]) );
	ao221_4 U293 ( .x(n94), .a(n102), .b(A[26]), .c(n102), .d(n109), .e(n108) );
	inv_2 U294 ( .x(n95), .a(n356) );
	nand2i_0 U295 ( .x(n356), .a(B[20]), .b(A[20]) );
	nand2i_2 U296 ( .x(n297), .a(n134), .b(n210) );
	nand2i_0 U297 ( .x(n111), .a(B[0]), .b(A[0]) );
	exnor2_1 U298 ( .x(n273), .a(A[18]), .b(B[18]) );
	nor2_0 U299 ( .x(n120), .a(n54), .b(n121) );
	nor2_0 U30 ( .x(n177), .a(n178), .b(n179) );
	nand2_2 U300 ( .x(n260), .a(n98), .b(n244) );
	inv_0 U301 ( .x(n250), .a(n98) );
	inv_10 U302 ( .x(n266), .a(n364) );
	nand4i_3 U303 ( .x(n268), .a(n148), .b(n338), .c(n339), .d(n340) );
	inv_0 U304 ( .x(n103), .a(n268) );
	inv_1 U305 ( .x(n104), .a(n103) );
	nand2i_4 U306 ( .x(n338), .a(n298), .b(n93) );
	exor2_1 U307 ( .x(DIFF[23]), .a(n104), .b(n269) );
	inv_2 U308 ( .x(n105), .a(n220) );
	exor2_1 U309 ( .x(n220), .a(A[31]), .b(B[31]) );
	exor2_1 U31 ( .x(DIFF[7]), .a(n215), .b(n122) );
	exor2_1 U310 ( .x(DIFF[16]), .a(n86), .b(n167) );
	aoi21_1 U311 ( .x(n199), .a(n86), .b(n200), .c(n311) );
	aoi21_1 U312 ( .x(n195), .a(n196), .b(n86), .c(n198) );
	aoi22_1 U313 ( .x(n203), .a(n204), .b(n205), .c(n206), .d(n86) );
	aoi21_1 U314 ( .x(n209), .a(n210), .b(n86), .c(n207) );
	inv_0 U315 ( .x(n335), .a(n258) );
	exnor2_1 U316 ( .x(DIFF[26]), .a(n264), .b(n265) );
	oai221_1 U317 ( .x(n223), .a(B[26]), .b(n264), .c(n264), .d(n238), .e(n343) );
	ao221_4 U319 ( .x(n212), .a(n101), .b(A[26]), .c(n101), .d(n109), .e(n108) );
	oai21_1 U32 ( .x(n215), .a(n127), .b(n327), .c(n319) );
	inv_2 U320 ( .x(n108), .a(n343) );
	inv_0 U321 ( .x(n109), .a(B[26]) );
	nand2i_0 U322 ( .x(n343), .a(B[26]), .b(A[26]) );
	inv_0 U323 ( .x(n238), .a(A[26]) );
	aoi21_3 U324 ( .x(n135), .a(n136), .b(n137), .c(n138) );
	exor2_3 U325 ( .x(DIFF[15]), .a(n227), .b(n169) );
	nand2_5 U326 ( .x(n253), .a(n254), .b(n78) );
	nand3i_3 U327 ( .x(n286), .a(n133), .b(n287), .c(n288) );
	nor2i_3 U328 ( .x(n305), .a(n306), .b(n211) );
	nor2i_3 U329 ( .x(n307), .a(A[29]), .b(n211) );
	inv_0 U33 ( .x(n127), .a(n236) );
	ao21_4 U330 ( .x(n227), .a(n228), .b(n248), .c(n173) );
	oai21_4 U331 ( .x(n137), .a(n126), .b(n124), .c(n235) );
	nand3i_3 U332 ( .x(n317), .a(n155), .b(n288), .c(n287) );
	nand2i_4 U333 ( .x(n328), .a(B[19]), .b(A[19]) );
	nand2i_4 U334 ( .x(n341), .a(B[23]), .b(A[23]) );
	nand2i_4 U337 ( .x(n339), .a(n300), .b(n357) );
	inv_5 U338 ( .x(n361), .a(n256) );
	oai21_4 U339 ( .x(n332), .a(n311), .b(n360), .c(n361) );
	inv_2 U34 ( .x(n327), .a(n216) );
	nand2i_4 U340 ( .x(n362), .a(n201), .b(n331) );
	nand2i_4 U341 ( .x(n363), .a(n149), .b(n268) );
	nand2_5 U342 ( .x(n364), .a(n363), .b(n341) );
	nand2_4 U344 ( .x(n340), .a(n337), .b(n299) );
	nand2i_6 U345 ( .x(n213), .a(A[27]), .b(B[27]) );
	nand2i_6 U346 ( .x(n249), .a(B[12]), .b(A[12]) );
	nand2i_5 U347 ( .x(n358), .a(n239), .b(n303) );
	aoi21_4 U348 ( .x(n301), .a(n302), .b(n303), .c(n304) );
	nand2i_6 U349 ( .x(n344), .a(B[27]), .b(A[27]) );
	nor2_1 U35 ( .x(n122), .a(n123), .b(n124) );
	nor2i_5 U350 ( .x(n114), .a(n115), .b(n116) );
	nand3i_1 U351 ( .x(n262), .a(n347), .b(n348), .c(n349) );
	nand3i_2 U352 ( .x(n351), .a(n308), .b(n348), .c(n349) );
	aoai211_3 U353 ( .x(n349), .a(n212), .b(n213), .c(n188), .d(n307) );
	or3i_5 U354 ( .x(n293), .a(n336), .b(n139), .c(n285) );
	nand4i_1 U355 ( .x(n350), .a(n87), .b(n349), .c(n348), .d(n309) );
	aoai211_3 U356 ( .x(n348), .a(n213), .b(n94), .c(n150), .d(n305) );
	nand2i_5 U357 ( .x(n316), .a(n232), .b(n277) );
	inv_0 U358 ( .x(n187), .a(n232) );
	nand2i_3 U359 ( .x(n232), .a(B[1]), .b(A[1]) );
	inv_2 U36 ( .x(n123), .a(n235) );
	inv_3 U360 ( .x(n100), .a(B[8]) );
	nand2i_2 U361 ( .x(n245), .a(A[8]), .b(B[8]) );
	inv_3 U362 ( .x(n58), .a(n313) );
	nand2i_3 U363 ( .x(n313), .a(B[10]), .b(A[10]) );
	nand2i_4 U364 ( .x(n197), .a(n295), .b(n292) );
	nand3i_5 U365 ( .x(n233), .a(n365), .b(n235), .c(n236) );
	inv_2 U366 ( .x(n365), .a(n234) );
	nand2i_3 U367 ( .x(n236), .a(A[6]), .b(B[6]) );
	nand2i_2 U368 ( .x(n235), .a(A[7]), .b(B[7]) );
	nand2_0 U369 ( .x(n141), .a(n83), .b(A[13]) );
	nand2_0 U37 ( .x(DIFF[0]), .a(n110), .b(n111) );
	inv_5 U370 ( .x(n83), .a(B[13]) );
	nand2i_2 U371 ( .x(n234), .a(A[5]), .b(B[5]) );
	inv_3 U372 ( .x(n85), .a(B[14]) );
	nand2i_4 U373 ( .x(n294), .a(A[15]), .b(B[15]) );
	nand2i_2 U374 ( .x(n319), .a(B[6]), .b(A[6]) );
	nor2i_0 U375 ( .x(n149), .a(B[23]), .b(A[23]) );
	inv_3 U376 ( .x(n67), .a(B[10]) );
	inv_5 U377 ( .x(n194), .a(B[18]) );
	nand2i_2 U378 ( .x(n252), .a(A[18]), .b(B[18]) );
	inv_0 U38 ( .x(n276), .a(n110) );
	nand2i_2 U39 ( .x(n243), .a(A[11]), .b(B[11]) );
	nor2i_1 U40 ( .x(n180), .a(n181), .b(n182) );
	oai21_1 U41 ( .x(n230), .a(n184), .b(n354), .c(n56) );
	inv_0 U42 ( .x(n89), .a(B[19]) );
	nor2i_1 U43 ( .x(n207), .a(n202), .b(n208) );
	nor2_0 U44 ( .x(n172), .a(n140), .b(n173) );
	inv_2 U45 ( .x(n140), .a(n248) );
	inv_2 U47 ( .x(n176), .a(n141) );
	or2_6 U48 ( .x(n247), .a(A[13]), .b(n83) );
	nor2_1 U49 ( .x(n174), .a(n82), .b(n176) );
	inv_2 U50 ( .x(n178), .a(n249) );
	oai21_1 U51 ( .x(n229), .a(n51), .b(n61), .c(n335) );
	inv_2 U52 ( .x(n353), .a(n229) );
	nand2i_2 U53 ( .x(n334), .a(A[12]), .b(B[12]) );
	oa21_2 U54 ( .x(n50), .a(n179), .b(n353), .c(n249) );
	nor2_1 U55 ( .x(n183), .a(n55), .b(n184) );
	inv_2 U56 ( .x(n354), .a(n231) );
	oai21_1 U57 ( .x(n231), .a(n324), .b(n119), .c(n325) );
	inv_0 U58 ( .x(n113), .a(n93) );
	nor2i_0 U59 ( .x(n112), .a(A[21]), .b(n113) );
	inv_0 U6 ( .x(n182), .a(n243) );
	inv_4 U60 ( .x(n96), .a(n362) );
	inv_2 U61 ( .x(n145), .a(B[21]) );
	nor2i_1 U62 ( .x(n144), .a(n145), .b(n113) );
	inv_2 U63 ( .x(n130), .a(n62) );
	nor2_1 U64 ( .x(n128), .a(n129), .b(n130) );
	oai21_1 U65 ( .x(n217), .a(n218), .b(n133), .c(n321) );
	nand2i_2 U66 ( .x(n318), .a(n114), .b(n317) );
	inv_2 U67 ( .x(n326), .a(n217) );
	inv_2 U68 ( .x(n166), .a(n314) );
	nor2_1 U69 ( .x(n206), .a(n251), .b(n166) );
	nand3_1 U7 ( .x(n116), .a(n277), .b(n110), .c(n278) );
	nand2i_0 U70 ( .x(n205), .a(n194), .b(n310) );
	nand2i_3 U72 ( .x(n330), .a(B[16]), .b(A[16]) );
	aoai211_1 U73 ( .x(n204), .a(n329), .b(n330), .c(n256), .d(n255) );
	nor2_1 U74 ( .x(n131), .a(n132), .b(n133) );
	inv_2 U75 ( .x(n132), .a(n321) );
	inv_2 U76 ( .x(n133), .a(n291) );
	nor2_1 U77 ( .x(n196), .a(n168), .b(n166) );
	nor2_1 U78 ( .x(n188), .a(n151), .b(n152) );
	inv_0 U79 ( .x(n306), .a(B[29]) );
	nand2_2 U8 ( .x(n323), .a(n322), .b(n321) );
	nor2_1 U80 ( .x(n150), .a(n151), .b(n152) );
	nand4_1 U81 ( .x(n136), .a(n62), .b(n235), .c(n323), .d(n236) );
	inv_2 U82 ( .x(n282), .a(n136) );
	inv_2 U83 ( .x(n124), .a(n320) );
	inv_2 U84 ( .x(n126), .a(n319) );
	nor2i_1 U85 ( .x(n281), .a(n137), .b(n282) );
	nand2i_2 U87 ( .x(n279), .a(n133), .b(n280) );
	inv_2 U88 ( .x(n151), .a(n345) );
	inv_2 U89 ( .x(n152), .a(n346) );
	nand2i_0 U9 ( .x(n320), .a(B[7]), .b(A[7]) );
	nand2i_2 U90 ( .x(n345), .a(n237), .b(n344) );
	nor2i_0 U91 ( .x(n189), .a(B[30]), .b(A[30]) );
	nand2i_2 U92 ( .x(n110), .a(A[0]), .b(B[0]) );
	aoi21_1 U93 ( .x(n185), .a(B[1]), .b(n186), .c(n187) );
	nand2i_2 U95 ( .x(n244), .a(A[9]), .b(B[9]) );
	inv_2 U96 ( .x(n119), .a(n244) );
	nor2_1 U97 ( .x(n117), .a(n118), .b(n119) );
	inv_2 U98 ( .x(n324), .a(n214) );
	inv_0 U99 ( .x(n99), .a(A[8]) );

endmodule


module EX_DW01_add_32_2_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire ___cell__39170_net140184, ___cell__39170_net140185, ___cell__39170_net140192,
	___cell__39170_net140193, ___cell__39170_net140197, ___cell__39170_net140199,
	___cell__39170_net140209, ___cell__39170_net140210, ___cell__39170_net140213,
	___cell__39170_net140214, ___cell__39170_net140218, ___cell__39170_net140223,
	___cell__39170_net140231, ___cell__39170_net140232, ___cell__39170_net140233,
	___cell__39170_net140235, ___cell__39170_net140236, ___cell__39170_net140238,
	___cell__39170_net140239, ___cell__39170_net140241, ___cell__39170_net140242,
	___cell__39170_net140244, ___cell__39170_net140246, ___cell__39170_net140249,
	___cell__39170_net140250, ___cell__39170_net140251, ___cell__39170_net140255,
	___cell__39170_net140256, ___cell__39170_net140257, ___cell__39170_net140258,
	___cell__39170_net140259, ___cell__39170_net140264, ___cell__39170_net140266,
	___cell__39170_net140267, ___cell__39170_net140268, ___cell__39170_net140269,
	___cell__39170_net140270, ___cell__39170_net140273, ___cell__39170_net140274,
	___cell__39170_net140276, ___cell__39170_net140277, ___cell__39170_net140278,
	___cell__39170_net140279, ___cell__39170_net140282, ___cell__39170_net140283,
	___cell__39170_net140284, ___cell__39170_net140285, ___cell__39170_net140286,
	___cell__39170_net140287, ___cell__39170_net140288, ___cell__39170_net140292,
	___cell__39170_net140305, ___cell__39170_net140307, ___cell__39170_net140309,
	___cell__39170_net140310, ___cell__39170_net140311, ___cell__39170_net140313,
	___cell__39170_net140316, ___cell__39170_net140317, ___cell__39170_net140319,
	___cell__39170_net140320, ___cell__39170_net140321, ___cell__39170_net140327,
	___cell__39170_net140337, ___cell__39170_net140341, ___cell__39170_net140351,
	___cell__39170_net140355, ___cell__39170_net140357, ___cell__39170_net140386,
	___cell__39170_net140392, ___cell__39170_net140395, ___cell__39170_net140396,
	___cell__39170_net140397, ___cell__39170_net140398, ___cell__39170_net140401,
	___cell__39170_net140410, ___cell__39170_net140411, ___cell__39170_net140412,
	___cell__39170_net140416, ___cell__39170_net140418, ___cell__39170_net140422,
	___cell__39170_net140424, ___cell__39170_net140427, ___cell__39170_net140444,
	___cell__39170_net140445, ___cell__39170_net140447, ___cell__39170_net140448,
	___cell__39170_net140451, ___cell__39170_net140452, ___cell__39170_net140455,
	___cell__39170_net140460, ___cell__39170_net140461, ___cell__39170_net140463,
	___cell__39170_net140464, ___cell__39170_net140471, ___cell__39170_net140476,
	___cell__39170_net140482, ___cell__39170_net140484, ___cell__39170_net140485,
	___cell__39170_net140490, ___cell__39170_net140495, ___cell__39170_net140499,
	___cell__39170_net140502, ___cell__39170_net140504, ___cell__39170_net140513,
	___cell__39170_net140514, ___cell__39170_net140525, ___cell__39170_net140528,
	___cell__39170_net140529, ___cell__39170_net140536, ___cell__39170_net140537,
	___cell__39170_net140541, ___cell__39170_net140546, ___cell__39170_net140560,
	___cell__39170_net140561, ___cell__39170_net140566, n100, n101, n102,
	n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
	n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
	n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
	n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
	n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
	n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173, n174,
	n175, n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
	n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
	n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
	n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
	n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233, n234,
	n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
	n247, n248, n249, n250, n251, n252, n49, n50, n51, n52, n53, n54, n55,
	n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
	n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
	n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
	n98, n99, net121836, net150005, net150142, net150555, net150690, net150837,
	net151030, net151031, net151032, net151417, net151951, net151953, net152445,
	net152474, net155899, net155900, net156215, net156380;


	inv_4 U10 ( .x(___cell__39170_net140238), .a(___cell__39170_net140310) );
	nor2i_1 U100 ( .x(n224), .a(n203), .b(n216) );
	inv_0 U101 ( .x(n203), .a(A[21]) );
	inv_0 U102 ( .x(n205), .a(B[20]) );
	exnor2_1 U103 ( .x(n223), .a(n216), .b(n203) );
	exor2_1 U104 ( .x(n180), .a(A[23]), .b(B[23]) );
	inv_2 U105 ( .x(___cell__39170_net140214), .a(___cell__39170_net140460) );
	inv_2 U106 ( .x(n202), .a(A[24]) );
	inv_2 U107 ( .x(n104), .a(A[23]) );
	nand2_2 U108 ( .x(___cell__39170_net140251), .a(B[23]), .b(A[23]) );
	exor2_1 U109 ( .x(___cell__39170_net140286), .a(B[25]), .b(A[25]) );
	inv_5 U11 ( .x(n98), .a(A[2]) );
	exor2_1 U110 ( .x(___cell__39170_net140285), .a(A[26]), .b(B[26]) );
	nand2_2 U111 ( .x(___cell__39170_net140357), .a(B[25]), .b(A[25]) );
	inv_2 U112 ( .x(___cell__39170_net140264), .a(___cell__39170_net140357) );
	inv_2 U113 ( .x(___cell__39170_net140355), .a(A[25]) );
	nand2i_2 U114 ( .x(n175), .a(B[25]), .b(___cell__39170_net140355) );
	exor2_1 U115 ( .x(SUM[3]), .a(___cell__39170_net140279), .b(___cell__39170_net140209) );
	nand3_1 U116 ( .x(___cell__39170_net140279), .a(___cell__39170_net140484),
		.b(n233), .c(n134) );
	nor2i_1 U117 ( .x(___cell__39170_net140209), .a(___cell__39170_net140210),
		.b(n121) );
	exnor2_1 U118 ( .x(SUM[2]), .a(n184), .b(n49) );
	nand2i_0 U119 ( .x(n184), .a(___cell__39170_net140238), .b(___cell__39170_net140316) );
	nand2i_4 U12 ( .x(___cell__39170_net140310), .a(B[2]), .b(n98) );
	inv_2 U120 ( .x(n245), .a(n247) );
	exor2_1 U121 ( .x(SUM[6]), .a(___cell__39170_net140273), .b(n144) );
	oai21_1 U122 ( .x(___cell__39170_net140273), .a(n120), .b(___cell__39170_net140502),
		.c(___cell__39170_net140193) );
	nor2i_0 U123 ( .x(n144), .a(n145), .b(n146) );
	inv_2 U124 ( .x(n168), .a(n150) );
	nor2i_0 U125 ( .x(n166), .a(n167), .b(n168) );
	inv_2 U126 ( .x(n70), .a(___cell__39170_net140246) );
	exor2_1 U127 ( .x(SUM[12]), .a(___cell__39170_net140199), .b(n166) );
	inv_0 U128 ( .x(n135), .a(n194) );
	nor2i_1 U129 ( .x(n141), .a(n142), .b(n135) );
	inv_2 U13 ( .x(___cell__39170_net140307), .a(B[0]) );
	inv_2 U130 ( .x(___cell__39170_net140504), .a(___cell__39170_net140273) );
	inv_0 U131 ( .x(n146), .a(n232) );
	oai21_1 U132 ( .x(n177), .a(n146), .b(___cell__39170_net140504), .c(n145) );
	exor2_1 U133 ( .x(SUM[7]), .a(n177), .b(n141) );
	inv_0 U134 ( .x(n56), .a(A[27]) );
	exor2_1 U135 ( .x(___cell__39170_net140284), .a(B[27]), .b(n58) );
	nor2i_1 U136 ( .x(SUM[0]), .a(n240), .b(n241) );
	exor2_1 U139 ( .x(SUM[20]), .a(net150837), .b(n183) );
	or3i_2 U14 ( .x(___cell__39170_net140309), .a(___cell__39170_net140310),
		.b(___cell__39170_net140305), .c(___cell__39170_net140307) );
	exor2_1 U140 ( .x(SUM[14]), .a(n191), .b(n163) );
	exnor2_1 U141 ( .x(SUM[13]), .a(n149), .b(n164) );
	aoi21_1 U142 ( .x(n149), .a(___cell__39170_net140199), .b(n150), .c(n151) );
	inv_2 U143 ( .x(n151), .a(n167) );
	nor2i_0 U144 ( .x(n164), .a(n165), .b(n91) );
	exor2_1 U146 ( .x(SUM[10]), .a(n193), .b(n169) );
	oai21_1 U147 ( .x(n193), .a(___cell__39170_net140269), .b(___cell__39170_net140185),
		.c(___cell__39170_net140184) );
	exor2_1 U149 ( .x(SUM[5]), .a(___cell__39170_net140274), .b(___cell__39170_net140192) );
	nand2i_1 U15 ( .x(n62), .a(___cell__39170_net140311), .b(___cell__39170_net140310) );
	oai21_1 U150 ( .x(___cell__39170_net140274), .a(___cell__39170_net140197),
		.b(n234), .c(n148) );
	nor2i_1 U151 ( .x(___cell__39170_net140192), .a(___cell__39170_net140193),
		.b(n120) );
	inv_2 U152 ( .x(___cell__39170_net140502), .a(___cell__39170_net140274) );
	exnor2_1 U153 ( .x(SUM[19]), .a(n157), .b(n185) );
	exor2_1 U154 ( .x(SUM[4]), .a(n178), .b(n147) );
	nand2i_2 U155 ( .x(n178), .a(___cell__39170_net140490), .b(___cell__39170_net140499) );
	inv_2 U156 ( .x(___cell__39170_net140490), .a(___cell__39170_net140210) );
	nor2i_1 U157 ( .x(n147), .a(n148), .b(___cell__39170_net140197) );
	inv_2 U158 ( .x(___cell__39170_net140197), .a(___cell__39170_net140321) );
	inv_2 U159 ( .x(n234), .a(n178) );
	nor2i_1 U16 ( .x(___cell__39170_net140445), .a(___cell__39170_net140444),
		.b(n62) );
	exor2_1 U161 ( .x(___cell__39170_net140282), .a(B[28]), .b(A[28]) );
	ao221_1 U162 ( .x(n179), .a(n50), .b(net151953), .c(n50), .d(n57), .e(net151951) );
	exor2_1 U163 ( .x(SUM[28]), .a(n179), .b(___cell__39170_net140282) );
	nor2i_1 U164 ( .x(n93), .a(n95), .b(n94) );
	inv_2 U165 ( .x(n94), .a(n231) );
	inv_5 U166 ( .x(net156380), .a(___cell__39170_net140267) );
	exnor2_1 U167 ( .x(SUM[1]), .a(n246), .b(n240) );
	exnor2_1 U168 ( .x(SUM[9]), .a(___cell__39170_net140269), .b(n140) );
	inv_2 U169 ( .x(___cell__39170_net140269), .a(___cell__39170_net140495) );
	inv_4 U17 ( .x(n125), .a(___cell__39170_net140319) );
	oai22_1 U170 ( .x(___cell__39170_net140495), .a(n112), .b(___cell__39170_net140341),
		.c(___cell__39170_net140395), .d(n93) );
	inv_2 U171 ( .x(n112), .a(B[8]) );
	inv_5 U172 ( .x(___cell__39170_net140341), .a(A[8]) );
	inv_5 U173 ( .x(___cell__39170_net140395), .a(___cell__39170_net140476) );
	nor2i_1 U174 ( .x(n140), .a(___cell__39170_net140184), .b(___cell__39170_net140185) );
	inv_2 U175 ( .x(___cell__39170_net140185), .a(___cell__39170_net140396) );
	inv_2 U176 ( .x(n236), .a(n191) );
	oai21_1 U177 ( .x(n189), .a(net152474), .b(n236), .c(___cell__39170_net140223) );
	exor2_1 U178 ( .x(SUM[15]), .a(n189), .b(n190) );
	exnor2_1 U179 ( .x(SUM[16]), .a(n188), .b(n160) );
	nor2i_3 U18 ( .x(___cell__39170_net140257), .a(___cell__39170_net140444),
		.b(___cell__39170_net140309) );
	nand2_2 U180 ( .x(SUM[21]), .a(n138), .b(n139) );
	nand2i_2 U181 ( .x(n139), .a(n154), .b(n216) );
	exnor2_1 U182 ( .x(SUM[23]), .a(___cell__39170_net140288), .b(n180) );
	exor2_1 U183 ( .x(SUM[24]), .a(___cell__39170_net140287), .b(n156) );
	or2_2 U184 ( .x(n49), .a(n243), .b(n245) );
	inv_2 U185 ( .x(n143), .a(n194) );
	nand2i_4 U186 ( .x(n194), .a(B[7]), .b(n196) );
	ao21_2 U187 ( .x(n50), .a(n97), .b(n51), .c(n106) );
	or2_2 U188 ( .x(n51), .a(n99), .b(n100) );
	nor2i_4 U189 ( .x(net152474), .a(n87), .b(A[14]) );
	nand2_0 U19 ( .x(n132), .a(A[19]), .b(B[19]) );
	nand2_2 U190 ( .x(n52), .a(n87), .b(n66) );
	nor2i_2 U191 ( .x(n61), .a(n89), .b(A[18]) );
	inv_3 U192 ( .x(___cell__39170_net140386), .a(B[15]) );
	inv_2 U193 ( .x(n53), .a(n54) );
	inv_2 U194 ( .x(n55), .a(n54) );
	inv_0 U195 ( .x(n57), .a(n56) );
	inv_0 U196 ( .x(n58), .a(n56) );
	inv_3 U197 ( .x(n124), .a(A[5]) );
	oai211_2 U198 ( .x(n220), .a(n188), .b(n72), .c(n217), .d(n250) );
	inv_2 U199 ( .x(n77), .a(n218) );
	nand2_2 U20 ( .x(___cell__39170_net140546), .a(A[29]), .b(B[29]) );
	inv_10 U200 ( .x(___cell__39170_net140320), .a(___cell__39170_net140317) );
	and3i_4 U201 ( .x(n82), .a(n214), .b(___cell__39170_net140242), .c(n52) );
	and3i_3 U202 ( .x(___cell__39170_net140244), .a(n79), .b(n88), .c(___cell__39170_net140242) );
	nand2i_3 U203 ( .x(___cell__39170_net140242), .a(A[15]), .b(___cell__39170_net140386) );
	or3i_3 U204 ( .x(n200), .a(___cell__39170_net140320), .b(___cell__39170_net140210),
		.c(n226) );
	nand2_2 U205 ( .x(n71), .a(n126), .b(n127) );
	inv_0 U206 ( .x(n59), .a(n238) );
	nand2i_2 U207 ( .x(n238), .a(B[16]), .b(n208) );
	inv_2 U208 ( .x(n162), .a(n238) );
	nand2_8 U209 ( .x(___cell__39170_net140317), .a(n232), .b(n194) );
	nand2i_2 U21 ( .x(___cell__39170_net140266), .a(A[29]), .b(n109) );
	or3i_3 U211 ( .x(___cell__39170_net140337), .a(___cell__39170_net140320),
		.b(n124), .c(___cell__39170_net140327) );
	inv_0 U212 ( .x(n210), .a(A[18]) );
	ao21_3 U214 ( .x(n63), .a(n145), .b(n142), .c(n143) );
	nand2_1 U215 ( .x(n142), .a(A[7]), .b(B[7]) );
	nand4_1 U216 ( .x(n198), .a(n199), .b(___cell__39170_net140337), .c(n200),
		.d(n63) );
	aoai211_1 U217 ( .x(___cell__39170_net140448), .a(n129), .b(n128), .c(n74),
		.d(n132) );
	inv_2 U218 ( .x(n64), .a(___cell__39170_net140471) );
	nand2_5 U219 ( .x(___cell__39170_net140258), .a(n88), .b(n82) );
	inv_4 U22 ( .x(n196), .a(A[7]) );
	inv_2 U220 ( .x(n66), .a(A[14]) );
	nor2i_0 U222 ( .x(___cell__39170_net140241), .a(___cell__39170_net140242),
		.b(n79) );
	aoi21_2 U223 ( .x(n79), .a(n65), .b(n133), .c(n130) );
	nand2_0 U224 ( .x(n148), .a(B[4]), .b(A[4]) );
	nand2i_2 U225 ( .x(___cell__39170_net140321), .a(A[4]), .b(n195) );
	nand2_0 U226 ( .x(n227), .a(B[4]), .b(A[4]) );
	inv_0 U227 ( .x(n209), .a(A[17]) );
	inv_6 U228 ( .x(___cell__39170_net140427), .a(___cell__39170_net140292) );
	inv_0 U229 ( .x(___cell__39170_net140327), .a(B[5]) );
	inv_2 U23 ( .x(n87), .a(B[14]) );
	aoai211_3 U230 ( .x(net150142), .a(___cell__39170_net140561), .b(___cell__39170_net140560),
		.c(___cell__39170_net140427), .d(___cell__39170_net140455) );
	or3i_2 U231 ( .x(n199), .a(___cell__39170_net140320), .b(n171), .c(n227) );
	exor2_1 U232 ( .x(n190), .a(A[15]), .b(B[15]) );
	nand2_0 U233 ( .x(n131), .a(A[15]), .b(B[15]) );
	ao211_5 U234 ( .x(___cell__39170_net140199), .a(n70), .b(n69), .c(n68),
		.d(n67) );
	inv_0 U235 ( .x(n67), .a(___cell__39170_net140514) );
	inv_0 U236 ( .x(n68), .a(___cell__39170_net140513) );
	inv_0 U237 ( .x(n69), .a(___cell__39170_net140259) );
	nor3_4 U238 ( .x(___cell__39170_net140246), .a(n172), .b(n173), .c(___cell__39170_net140249) );
	inv_4 U239 ( .x(n122), .a(n71) );
	inv_0 U24 ( .x(n155), .a(A[22]) );
	inv_0 U240 ( .x(n121), .a(n127) );
	inv_0 U241 ( .x(n120), .a(n126) );
	nand2i_2 U242 ( .x(n126), .a(B[5]), .b(n124) );
	nand2i_0 U243 ( .x(n72), .a(n162), .b(n212) );
	nand2i_4 U244 ( .x(n211), .a(n162), .b(n212) );
	nand2i_2 U245 ( .x(n212), .a(B[17]), .b(n209) );
	inv_6 U246 ( .x(n215), .a(A[11]) );
	nor2i_1 U248 ( .x(n114), .a(A[8]), .b(n112) );
	inv_0 U249 ( .x(n73), .a(___cell__39170_net140311) );
	inv_2 U25 ( .x(n153), .a(B[22]) );
	nor3_2 U250 ( .x(___cell__39170_net140451), .a(___cell__39170_net140448),
		.b(___cell__39170_net140244), .c(___cell__39170_net140256) );
	inv_0 U251 ( .x(___cell__39170_net140218), .a(n74) );
	inv_4 U252 ( .x(n197), .a(B[6]) );
	inv_2 U253 ( .x(n133), .a(net152474) );
	inv_2 U254 ( .x(n80), .a(___cell__39170_net140445) );
	inv_2 U255 ( .x(n81), .a(n172) );
	exnor2_5 U256 ( .x(SUM[30]), .a(n83), .b(n96) );
	inv_0 U257 ( .x(___cell__39170_net140401), .a(n82) );
	nand2i_2 U258 ( .x(n237), .a(___cell__39170_net140401), .b(___cell__39170_net140199) );
	nand2_5 U259 ( .x(___cell__39170_net140566), .a(n51), .b(n97) );
	aoi21_1 U26 ( .x(n152), .a(n153), .b(n154), .c(n155) );
	nand3_2 U260 ( .x(___cell__39170_net140292), .a(___cell__39170_net140451),
		.b(___cell__39170_net140452), .c(___cell__39170_net140525) );
	ao21_4 U261 ( .x(n83), .a(___cell__39170_net140267), .b(___cell__39170_net140266),
		.c(___cell__39170_net140268) );
	inv_2 U263 ( .x(n85), .a(B[13]) );
	inv_10 U264 ( .x(n86), .a(A[6]) );
	nand2i_2 U265 ( .x(___cell__39170_net140397), .a(B[10]), .b(n113) );
	nor2_6 U266 ( .x(n88), .a(___cell__39170_net140392), .b(n211) );
	nand4_1 U268 ( .x(___cell__39170_net140412), .a(___cell__39170_net140398),
		.b(___cell__39170_net140396), .c(n114), .d(n60) );
	inv_0 U269 ( .x(___cell__39170_net140236), .a(n60) );
	nand2_5 U27 ( .x(n207), .a(A[20]), .b(B[20]) );
	inv_2 U272 ( .x(n90), .a(n89) );
	aoai211_3 U274 ( .x(n108), .a(___cell__39170_net140561), .b(___cell__39170_net140560),
		.c(___cell__39170_net140427), .d(___cell__39170_net140455) );
	exnor2_3 U275 ( .x(SUM[31]), .a(___cell__39170_net140276), .b(net150005) );
	ao21_3 U276 ( .x(___cell__39170_net140525), .a(___cell__39170_net140514),
		.b(___cell__39170_net140513), .c(___cell__39170_net140258) );
	nor2i_1 U277 ( .x(n156), .a(___cell__39170_net140213), .b(___cell__39170_net140214) );
	inv_2 U278 ( .x(net150690), .a(net156215) );
	buf_2 U279 ( .x(net151417), .a(n97) );
	inv_2 U28 ( .x(n228), .a(n207) );
	inv_2 U280 ( .x(n208), .a(A[16]) );
	inv_2 U281 ( .x(___cell__39170_net140482), .a(___cell__39170_net140309) );
	inv_0 U282 ( .x(___cell__39170_net140270), .a(n93) );
	inv_0 U283 ( .x(n95), .a(n198) );
	nand2_0 U284 ( .x(___cell__39170_net140193), .a(B[5]), .b(A[5]) );
	nor2_0 U285 ( .x(n171), .a(B[5]), .b(A[5]) );
	oai22_1 U286 ( .x(n226), .a(A[4]), .b(B[4]), .c(B[5]), .d(A[5]) );
	inv_2 U287 ( .x(n96), .a(___cell__39170_net140278) );
	nand4i_3 U288 ( .x(n97), .a(___cell__39170_net140250), .b(___cell__39170_net140528),
		.c(___cell__39170_net140529), .d(___cell__39170_net140213) );
	nand2_1 U289 ( .x(n217), .a(B[17]), .b(A[17]) );
	nand2_2 U29 ( .x(___cell__39170_net140561), .a(n229), .b(B[20]) );
	nand2i_4 U290 ( .x(___cell__39170_net140528), .a(___cell__39170_net140461),
		.b(n108) );
	exor3_1 U291 ( .x(SUM[29]), .a(A[29]), .b(B[29]), .c(___cell__39170_net140267) );
	aoai211_1 U292 ( .x(___cell__39170_net140287), .a(n104), .b(___cell__39170_net140416),
		.c(___cell__39170_net140288), .d(___cell__39170_net140251) );
	inv_2 U293 ( .x(___cell__39170_net140416), .a(B[23]) );
	inv_0 U294 ( .x(___cell__39170_net140288), .a(n108) );
	inv_3 U295 ( .x(___cell__39170_net140305), .a(A[0]) );
	nand2i_2 U296 ( .x(___cell__39170_net140313), .a(___cell__39170_net140311),
		.b(___cell__39170_net140310) );
	nand2_2 U297 ( .x(___cell__39170_net140316), .a(B[2]), .b(A[2]) );
	inv_0 U298 ( .x(net155900), .a(B[1]) );
	nand2i_6 U299 ( .x(___cell__39170_net140283), .a(n106), .b(___cell__39170_net140566) );
	nand2i_2 U30 ( .x(n105), .a(n104), .b(___cell__39170_net140460) );
	nand2i_4 U300 ( .x(___cell__39170_net140536), .a(___cell__39170_net140464),
		.b(___cell__39170_net140283) );
	oai22_3 U301 ( .x(n106), .a(n101), .b(___cell__39170_net140357), .c(___cell__39170_net140351),
		.d(n102) );
	nand2i_4 U302 ( .x(___cell__39170_net140529), .a(n105), .b(net150142) );
	inv_0 U303 ( .x(net156215), .a(___cell__39170_net140427) );
	nand3i_3 U304 ( .x(___cell__39170_net140410), .a(___cell__39170_net140411),
		.b(___cell__39170_net140412), .c(n103) );
	aoi31_1 U305 ( .x(n103), .a(n60), .b(___cell__39170_net140398), .c(___cell__39170_net140447),
		.d(___cell__39170_net140239) );
	ao221_4 U306 ( .x(___cell__39170_net140276), .a(n111), .b(net151032), .c(n111),
		.d(net151031), .e(net151030) );
	inv_2 U307 ( .x(net151030), .a(___cell__39170_net140541) );
	nand2_0 U308 ( .x(___cell__39170_net140541), .a(A[30]), .b(B[30]) );
	inv_2 U309 ( .x(net151031), .a(___cell__39170_net140424) );
	nand2i_2 U31 ( .x(___cell__39170_net140461), .a(___cell__39170_net140416),
		.b(___cell__39170_net140460) );
	inv_2 U310 ( .x(___cell__39170_net140424), .a(A[30]) );
	inv_2 U311 ( .x(net151032), .a(___cell__39170_net140422) );
	inv_0 U312 ( .x(___cell__39170_net140422), .a(B[30]) );
	aoai211_4 U313 ( .x(n111), .a(n110), .b(n109), .c(net156380), .d(___cell__39170_net140546) );
	inv_6 U314 ( .x(n109), .a(B[29]) );
	exor2_1 U315 ( .x(___cell__39170_net140278), .a(B[30]), .b(A[30]) );
	nor2_2 U316 ( .x(___cell__39170_net140239), .a(___cell__39170_net140233),
		.b(___cell__39170_net140235) );
	nand4i_5 U317 ( .x(___cell__39170_net140267), .a(n115), .b(___cell__39170_net140536),
		.c(___cell__39170_net140537), .d(n119) );
	inv_0 U318 ( .x(___cell__39170_net140418), .a(B[27]) );
	nand2_0 U319 ( .x(___cell__39170_net140255), .a(n57), .b(B[27]) );
	nor2_1 U32 ( .x(___cell__39170_net140250), .a(___cell__39170_net140214),
		.b(___cell__39170_net140251) );
	inv_0 U320 ( .x(net150555), .a(n125) );
	nand3_4 U321 ( .x(___cell__39170_net140319), .a(___cell__39170_net140320),
		.b(___cell__39170_net140321), .c(n122) );
	inv_2 U322 ( .x(net151951), .a(___cell__39170_net140255) );
	nand2_2 U323 ( .x(n130), .a(n131), .b(___cell__39170_net140223) );
	inv_10 U324 ( .x(n128), .a(B[19]) );
	inv_2 U325 ( .x(net150005), .a(___cell__39170_net140277) );
	exor2_1 U326 ( .x(___cell__39170_net140277), .a(B[31]), .b(A[31]) );
	aoi21_1 U327 ( .x(n174), .a(n175), .b(net151417), .c(___cell__39170_net140264) );
	exor2_1 U328 ( .x(SUM[25]), .a(net151417), .b(___cell__39170_net140286) );
	nor2_0 U329 ( .x(n134), .a(net152445), .b(n170) );
	and4i_3 U33 ( .x(n170), .a(___cell__39170_net140238), .b(A[0]), .c(B[0]),
		.d(A[1]) );
	nand2_0 U330 ( .x(n240), .a(A[0]), .b(B[0]) );
	and3i_1 U331 ( .x(n243), .a(n244), .b(B[0]), .c(A[0]) );
	nor2_0 U332 ( .x(n241), .a(B[0]), .b(A[0]) );
	or2_6 U333 ( .x(n172), .a(n170), .b(net152445) );
	nand2_0 U334 ( .x(n219), .a(B[18]), .b(A[18]) );
	nor2i_2 U335 ( .x(n225), .a(A[18]), .b(n220) );
	inv_2 U336 ( .x(net151953), .a(___cell__39170_net140418) );
	exor2_1 U337 ( .x(SUM[27]), .a(n50), .b(___cell__39170_net140284) );
	nand2i_2 U338 ( .x(___cell__39170_net140460), .a(B[24]), .b(n202) );
	nand2_0 U339 ( .x(___cell__39170_net140213), .a(A[24]), .b(B[24]) );
	inv_1 U34 ( .x(___cell__39170_net140311), .a(A[1]) );
	exor2_1 U340 ( .x(n187), .a(B[17]), .b(A[17]) );
	ao21_1 U341 ( .x(n176), .a(A[8]), .b(B[8]), .c(___cell__39170_net140395) );
	inv_0 U342 ( .x(net150837), .a(net150690) );
	inv_3 U343 ( .x(n201), .a(B[9]) );
	nand2_3 U344 ( .x(___cell__39170_net140184), .a(B[9]), .b(A[9]) );
	exnor2_1 U345 ( .x(SUM[8]), .a(___cell__39170_net140270), .b(n176) );
	oai22_1 U346 ( .x(n206), .a(B[21]), .b(A[21]), .c(A[22]), .d(B[22]) );
	nand2_4 U347 ( .x(n154), .a(B[21]), .b(A[21]) );
	mux2i_1 U348 ( .x(n138), .d0(n223), .sl(B[21]), .d1(n224) );
	inv_0 U349 ( .x(n204), .a(B[21]) );
	nor2_1 U35 ( .x(n244), .a(net121836), .b(n73) );
	oai211_1 U350 ( .x(n218), .a(A[17]), .b(B[17]), .c(A[16]), .d(B[16]) );
	nand2_0 U351 ( .x(n161), .a(A[16]), .b(B[16]) );
	nor2i_0 U352 ( .x(n169), .a(n64), .b(___cell__39170_net140236) );
	inv_0 U353 ( .x(___cell__39170_net140471), .a(___cell__39170_net140235) );
	inv_3 U355 ( .x(n213), .a(B[12]) );
	nand2_0 U356 ( .x(___cell__39170_net140235), .a(A[10]), .b(B[10]) );
	exnor2_3 U357 ( .x(SUM[26]), .a(n174), .b(___cell__39170_net140285) );
	nand2i_4 U358 ( .x(n214), .a(n168), .b(n84) );
	exnor2_3 U359 ( .x(n221), .a(n222), .b(n210) );
	nand2i_4 U36 ( .x(___cell__39170_net140259), .a(n92), .b(n125) );
	aoi221_4 U360 ( .x(___cell__39170_net140455), .a(n228), .b(n229), .c(B[22]),
		.d(n230), .e(n152) );
	nand2i_4 U361 ( .x(___cell__39170_net140476), .a(B[8]), .b(___cell__39170_net140341) );
	mux2i_3 U363 ( .x(n136), .d0(n225), .sl(n90), .d1(n221) );
	nand2_3 U364 ( .x(SUM[18]), .a(n136), .b(n137) );
	aoai211_5 U365 ( .x(n216), .a(n205), .b(n54), .c(net150690), .d(n207) );
	nand2i_6 U366 ( .x(___cell__39170_net140398), .a(B[11]), .b(n215) );
	nand2_8 U367 ( .x(___cell__39170_net140560), .a(n229), .b(n53) );
	inv_6 U368 ( .x(n229), .a(n206) );
	inv_10 U369 ( .x(n195), .a(B[4]) );
	inv_2 U37 ( .x(___cell__39170_net140444), .a(net155899) );
	inv_2 U370 ( .x(net121836), .a(net155900) );
	or2_2 U371 ( .x(n137), .a(n76), .b(n222) );
	inv_3 U372 ( .x(n222), .a(n220) );
	exnor2_1 U373 ( .x(SUM[22]), .a(n181), .b(n248) );
	inv_2 U374 ( .x(n248), .a(n182) );
	aoai211_2 U375 ( .x(n181), .a(n204), .b(n203), .c(n239), .d(n154) );
	ao211_4 U376 ( .x(___cell__39170_net140452), .a(n80), .b(n81), .c(___cell__39170_net140258),
		.d(___cell__39170_net140259) );
	exnor2_3 U377 ( .x(SUM[11]), .a(n249), .b(___cell__39170_net140231) );
	inv_3 U378 ( .x(n249), .a(n192) );
	ao21_2 U379 ( .x(n192), .a(n193), .b(n60), .c(___cell__39170_net140471) );
	inv_2 U38 ( .x(___cell__39170_net140485), .a(___cell__39170_net140313) );
	nor2i_0 U380 ( .x(___cell__39170_net140231), .a(___cell__39170_net140232),
		.b(___cell__39170_net140233) );
	inv_2 U381 ( .x(n113), .a(A[10]) );
	ao21_3 U382 ( .x(___cell__39170_net140392), .a(n128), .b(n129), .c(n61) );
	inv_4 U383 ( .x(n129), .a(A[19]) );
	nand4i_2 U384 ( .x(n92), .a(___cell__39170_net140395), .b(___cell__39170_net140396),
		.c(n60), .d(___cell__39170_net140398) );
	buf_8 U385 ( .x(n60), .a(___cell__39170_net140397) );
	nor3i_4 U386 ( .x(___cell__39170_net140256), .a(___cell__39170_net140257),
		.b(___cell__39170_net140259), .c(___cell__39170_net140258) );
	inv_0 U387 ( .x(n250), .a(n77) );
	oaoi211_2 U388 ( .x(n74), .a(n78), .b(n77), .c(n76), .d(n75) );
	ao21_4 U389 ( .x(n65), .a(n84), .b(n151), .c(n251) );
	nand2_2 U39 ( .x(___cell__39170_net140484), .a(___cell__39170_net140485),
		.b(___cell__39170_net140444) );
	inv_0 U390 ( .x(n91), .a(n84) );
	inv_0 U391 ( .x(n165), .a(n251) );
	nor2i_1 U392 ( .x(n251), .a(B[13]), .b(n252) );
	nand2i_2 U393 ( .x(n84), .a(A[13]), .b(n85) );
	inv_1 U394 ( .x(n252), .a(A[13]) );
	inv_2 U40 ( .x(___cell__39170_net140249), .a(___cell__39170_net140484) );
	inv_2 U41 ( .x(net155899), .a(B[1]) );
	nand2i_2 U42 ( .x(n233), .a(net155899), .b(___cell__39170_net140482) );
	inv_2 U43 ( .x(n173), .a(n233) );
	inv_2 U44 ( .x(net152445), .a(___cell__39170_net140316) );
	nand2i_5 U45 ( .x(n232), .a(A[6]), .b(n197) );
	or2_5 U46 ( .x(n145), .a(n86), .b(n197) );
	inv_2 U47 ( .x(___cell__39170_net140351), .a(B[26]) );
	inv_2 U48 ( .x(n102), .a(A[26]) );
	nand2i_2 U49 ( .x(n107), .a(B[26]), .b(n102) );
	nor2i_1 U50 ( .x(n99), .a(B[25]), .b(n101) );
	inv_2 U51 ( .x(n101), .a(n107) );
	nor2i_0 U52 ( .x(n100), .a(A[25]), .b(n101) );
	inv_2 U53 ( .x(___cell__39170_net140233), .a(___cell__39170_net140398) );
	inv_2 U54 ( .x(___cell__39170_net140411), .a(___cell__39170_net140232) );
	nand2_0 U55 ( .x(___cell__39170_net140232), .a(A[11]), .b(B[11]) );
	exor2_1 U56 ( .x(n183), .a(n55), .b(B[20]) );
	inv_2 U57 ( .x(n54), .a(A[20]) );
	nor2i_1 U58 ( .x(n163), .a(___cell__39170_net140223), .b(net152474) );
	nand2_1 U59 ( .x(n167), .a(A[12]), .b(B[12]) );
	nand2i_4 U6 ( .x(___cell__39170_net140513), .a(n92), .b(n198) );
	nand2i_5 U60 ( .x(n150), .a(A[12]), .b(n213) );
	exor2_1 U61 ( .x(n182), .a(A[22]), .b(B[22]) );
	exor2_1 U63 ( .x(n185), .a(A[19]), .b(B[19]) );
	aoi21_1 U64 ( .x(n157), .a(n158), .b(n159), .c(___cell__39170_net140218) );
	nor2i_1 U65 ( .x(n158), .a(n76), .b(n72) );
	inv_2 U66 ( .x(n76), .a(n61) );
	inv_2 U68 ( .x(n78), .a(n217) );
	inv_2 U69 ( .x(n75), .a(n219) );
	inv_5 U7 ( .x(___cell__39170_net140514), .a(___cell__39170_net140410) );
	nand2_1 U70 ( .x(___cell__39170_net140210), .a(A[3]), .b(B[3]) );
	nand2i_2 U71 ( .x(___cell__39170_net140499), .a(n121), .b(___cell__39170_net140279) );
	nand2i_2 U72 ( .x(n127), .a(B[3]), .b(n123) );
	inv_2 U73 ( .x(n123), .a(A[3]) );
	inv_2 U74 ( .x(n188), .a(n159) );
	nand2i_2 U75 ( .x(n231), .a(net150555), .b(___cell__39170_net140279) );
	nand2_2 U76 ( .x(n119), .a(B[28]), .b(A[28]) );
	nand2i_4 U77 ( .x(___cell__39170_net140537), .a(___cell__39170_net140463),
		.b(___cell__39170_net140283) );
	nand2i_2 U78 ( .x(___cell__39170_net140463), .a(n116), .b(B[27]) );
	nand2i_2 U79 ( .x(___cell__39170_net140464), .a(n116), .b(n58) );
	inv_7 U8 ( .x(n89), .a(B[18]) );
	inv_2 U80 ( .x(n117), .a(B[28]) );
	nand2i_2 U81 ( .x(n118), .a(A[28]), .b(n117) );
	inv_2 U82 ( .x(n116), .a(n118) );
	nor2_1 U83 ( .x(n115), .a(n116), .b(___cell__39170_net140255) );
	inv_2 U84 ( .x(___cell__39170_net140268), .a(___cell__39170_net140546) );
	inv_2 U85 ( .x(n110), .a(A[29]) );
	nor2_1 U86 ( .x(n242), .a(net121836), .b(n73) );
	nand2_2 U87 ( .x(n247), .a(n73), .b(net121836) );
	nor2i_1 U88 ( .x(n246), .a(n247), .b(n242) );
	nand2i_2 U89 ( .x(___cell__39170_net140396), .a(A[9]), .b(n201) );
	inv_2 U90 ( .x(___cell__39170_net140447), .a(___cell__39170_net140184) );
	nand2i_0 U91 ( .x(n235), .a(n214), .b(___cell__39170_net140199) );
	nand2i_2 U92 ( .x(n191), .a(n65), .b(n235) );
	nand2_1 U93 ( .x(___cell__39170_net140223), .a(A[14]), .b(B[14]) );
	nand2i_2 U94 ( .x(n159), .a(___cell__39170_net140241), .b(n237) );
	nor2i_1 U95 ( .x(n160), .a(n161), .b(n59) );
	exor2_1 U96 ( .x(SUM[17]), .a(n186), .b(n187) );
	oai21_1 U97 ( .x(n186), .a(n188), .b(n59), .c(n161) );
	inv_2 U98 ( .x(n230), .a(n154) );
	inv_2 U99 ( .x(n239), .a(n216) );

endmodule


module EX_DW01_add_32_0_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
	n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n268,
	n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
	n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
	n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
	n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
	n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328,
	n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
	n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
	n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
	n365, n366, n367, n368, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
	n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
	n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
	n87, n88, n89, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	inv_2 U10 ( .x(n119), .a(n301) );
	inv_2 U100 ( .x(n79), .a(n323) );
	mux2i_1 U101 ( .x(n109), .d0(n287), .sl(B[1]), .d1(n289) );
	nand2i_2 U102 ( .x(n191), .a(n115), .b(n332) );
	nor2i_0 U103 ( .x(n115), .a(A[8]), .b(n116) );
	nand2_2 U104 ( .x(n332), .a(n192), .b(n325) );
	inv_2 U105 ( .x(n333), .a(n191) );
	nor2i_1 U107 ( .x(n165), .a(n63), .b(n167) );
	inv_2 U108 ( .x(n280), .a(n139) );
	oai21_1 U109 ( .x(n279), .a(n167), .b(n280), .c(n63) );
	nand3_1 U11 ( .x(n272), .a(n185), .b(n301), .c(n302) );
	nand2_4 U110 ( .x(n93), .a(n95), .b(n248) );
	nand2i_2 U111 ( .x(n113), .a(n281), .b(n279) );
	exnor2_1 U112 ( .x(n285), .a(n286), .b(n95) );
	inv_2 U113 ( .x(n286), .a(n279) );
	inv_8 U114 ( .x(n95), .a(B[17]) );
	nor2i_1 U115 ( .x(n154), .a(n155), .b(n156) );
	nand2_2 U116 ( .x(n155), .a(B[21]), .b(A[21]) );
	inv_2 U117 ( .x(n246), .a(B[21]) );
	inv_2 U118 ( .x(n105), .a(n276) );
	inv_2 U119 ( .x(n106), .a(n253) );
	inv_1 U12 ( .x(n173), .a(n259) );
	inv_2 U120 ( .x(n158), .a(n260) );
	nand2i_2 U121 ( .x(n261), .a(n136), .b(n158) );
	inv_2 U122 ( .x(n252), .a(B[19]) );
	exor2_1 U123 ( .x(n206), .a(B[23]), .b(A[23]) );
	inv_0 U124 ( .x(n238), .a(A[24]) );
	inv_2 U125 ( .x(n235), .a(A[26]) );
	inv_2 U127 ( .x(n153), .a(n241) );
	inv_2 U128 ( .x(n236), .a(A[25]) );
	nand2i_2 U129 ( .x(n347), .a(B[25]), .b(n236) );
	inv_0 U13 ( .x(n170), .a(n257) );
	inv_3 U130 ( .x(n108), .a(n80) );
	exor2_1 U131 ( .x(SUM[3]), .a(n198), .b(n148) );
	exnor2_1 U132 ( .x(SUM[2]), .a(n209), .b(n51) );
	nand2i_2 U133 ( .x(n209), .a(n233), .b(n234) );
	exor2_1 U134 ( .x(SUM[6]), .a(n121), .b(n126) );
	nor2i_1 U135 ( .x(n174), .a(n175), .b(n176) );
	exor2_1 U136 ( .x(SUM[12]), .a(n216), .b(n174) );
	exnor2_1 U137 ( .x(SUM[7]), .a(n120), .b(n124) );
	aoi21_1 U138 ( .x(n120), .a(n121), .b(n122), .c(n123) );
	nor2i_1 U139 ( .x(n124), .a(n125), .b(n87) );
	nand2i_0 U14 ( .x(n259), .a(A[13]), .b(n270) );
	exnor2_1 U140 ( .x(SUM[27]), .a(n201), .b(n202) );
	exor2_1 U141 ( .x(SUM[11]), .a(n217), .b(n177) );
	exnor2_1 U142 ( .x(SUM[20]), .a(n157), .b(n208) );
	exor2_1 U143 ( .x(SUM[14]), .a(n214), .b(n168) );
	oai21_1 U144 ( .x(n214), .a(n173), .b(n353), .c(n172) );
	nor2i_1 U145 ( .x(n168), .a(n169), .b(n170) );
	inv_2 U146 ( .x(n354), .a(n214) );
	exor2_1 U147 ( .x(SUM[13]), .a(n215), .b(n171) );
	inv_2 U148 ( .x(n176), .a(n258) );
	nor2i_1 U149 ( .x(n171), .a(n172), .b(n173) );
	nand4i_1 U15 ( .x(n255), .a(n256), .b(n257), .c(n258), .d(n259) );
	inv_2 U150 ( .x(n353), .a(n215) );
	exor2_1 U151 ( .x(SUM[10]), .a(n218), .b(n180) );
	inv_2 U152 ( .x(n335), .a(n194) );
	nor2i_1 U153 ( .x(n129), .a(n130), .b(n131) );
	oai21_1 U154 ( .x(n194), .a(n134), .b(n334), .c(n133) );
	exor2_1 U155 ( .x(SUM[5]), .a(n194), .b(n129) );
	exnor2_1 U156 ( .x(SUM[19]), .a(n160), .b(n210) );
	exor2_1 U157 ( .x(SUM[4]), .a(n195), .b(n132) );
	oai21_1 U158 ( .x(n195), .a(n150), .b(n329), .c(n149) );
	inv_2 U159 ( .x(n150), .a(n326) );
	nand2_1 U16 ( .x(n118), .a(B[9]), .b(A[9]) );
	inv_2 U160 ( .x(n329), .a(n198) );
	nor2i_1 U161 ( .x(n132), .a(n133), .b(n134) );
	inv_2 U162 ( .x(n334), .a(n195) );
	exnor2_1 U163 ( .x(SUM[18]), .a(n162), .b(n211) );
	inv_2 U164 ( .x(n349), .a(n348) );
	exor2_1 U165 ( .x(n200), .a(B[28]), .b(n59) );
	inv_2 U166 ( .x(n317), .a(n325) );
	exnor2_1 U167 ( .x(SUM[8]), .a(n192), .b(n193) );
	exnor2_1 U168 ( .x(SUM[29]), .a(n283), .b(n284) );
	nand2_2 U169 ( .x(SUM[1]), .a(n109), .b(n53) );
	nand3_1 U17 ( .x(n356), .a(n259), .b(n257), .c(n339) );
	exor2_1 U170 ( .x(SUM[9]), .a(n191), .b(n117) );
	exor2_1 U171 ( .x(SUM[15]), .a(n212), .b(n213) );
	exor2_1 U172 ( .x(SUM[16]), .a(n139), .b(n165) );
	nand2_2 U173 ( .x(SUM[17]), .a(n112), .b(n113) );
	exnor2_1 U174 ( .x(SUM[21]), .a(n137), .b(n154) );
	inv_2 U175 ( .x(n358), .a(n242) );
	nand2i_2 U176 ( .x(n204), .a(n240), .b(n237) );
	inv_2 U177 ( .x(n232), .a(B[9]) );
	inv_2 U178 ( .x(n247), .a(B[16]) );
	inv_0 U179 ( .x(n116), .a(B[8]) );
	nand2i_2 U18 ( .x(n359), .a(n172), .b(n257) );
	inv_2 U180 ( .x(n318), .a(B[28]) );
	or2_2 U181 ( .x(n51), .a(n361), .b(n363) );
	inv_2 U182 ( .x(n290), .a(n87) );
	and2_3 U183 ( .x(n87), .a(n88), .b(n227) );
	aoi21_4 U184 ( .x(n52), .a(n296), .b(n302), .c(n189) );
	or2_2 U185 ( .x(n53), .a(n364), .b(n110) );
	inv_2 U186 ( .x(n156), .a(n337) );
	nand2i_2 U187 ( .x(n337), .a(A[21]), .b(n246) );
	nand2_2 U188 ( .x(n54), .a(n348), .b(n319) );
	nand2_2 U189 ( .x(n55), .a(n348), .b(n318) );
	oai22_3 U190 ( .x(n164), .a(n95), .b(n248), .c(n94), .d(n166) );
	ao21_4 U191 ( .x(n56), .a(n363), .b(n223), .c(n365) );
	inv_2 U192 ( .x(n363), .a(n364) );
	and4_3 U193 ( .x(n57), .a(n326), .b(n122), .c(n220), .d(n221) );
	inv_2 U194 ( .x(n273), .a(n77) );
	oa211_2 U195 ( .x(n77), .a(n239), .b(n242), .c(n274), .d(n152) );
	exor2_1 U196 ( .x(n213), .a(B[15]), .b(A[15]) );
	nand2i_2 U197 ( .x(n300), .a(B[15]), .b(n268) );
	nand2i_0 U198 ( .x(n346), .a(B[24]), .b(n238) );
	exor2_1 U199 ( .x(n205), .a(B[24]), .b(A[24]) );
	nor2i_3 U200 ( .x(n308), .a(A[30]), .b(n146) );
	inv_4 U201 ( .x(n146), .a(n352) );
	exnor2_1 U202 ( .x(SUM[23]), .a(n101), .b(n206) );
	aoi21_1 U203 ( .x(n157), .a(n158), .b(n139), .c(n103) );
	oai21_3 U204 ( .x(n143), .a(n156), .b(n104), .c(n155) );
	ao211_5 U205 ( .x(n295), .a(n133), .b(n130), .c(n128), .d(n131) );
	aoai211_4 U206 ( .x(n96), .a(n55), .b(n54), .c(n74), .d(n97) );
	inv_2 U207 ( .x(n59), .a(n319) );
	inv_2 U208 ( .x(n319), .a(A[28]) );
	nor3_2 U209 ( .x(n303), .a(n190), .b(n263), .c(n271) );
	nor2_0 U21 ( .x(n135), .a(A[19]), .b(B[19]) );
	aoi21_3 U210 ( .x(n190), .a(n58), .b(A[0]), .c(n84) );
	nand2i_2 U211 ( .x(n315), .a(n189), .b(n188) );
	ao21_1 U212 ( .x(n201), .a(n108), .b(n322), .c(n273) );
	nand2_0 U213 ( .x(n172), .a(B[13]), .b(A[13]) );
	oai22_2 U214 ( .x(n60), .a(n95), .b(n248), .c(n166), .d(n94) );
	inv_7 U215 ( .x(n94), .a(n93) );
	inv_2 U216 ( .x(n228), .a(A[5]) );
	nand2i_4 U217 ( .x(n321), .a(B[29]), .b(n96) );
	nor2i_0 U218 ( .x(n289), .a(n110), .b(A[1]) );
	nor2_0 U219 ( .x(n362), .a(B[1]), .b(A[1]) );
	inv_3 U22 ( .x(n92), .a(n60) );
	exnor2_1 U220 ( .x(n287), .a(A[1]), .b(n110) );
	nand2_2 U221 ( .x(n364), .a(B[1]), .b(A[1]) );
	inv_2 U222 ( .x(n73), .a(A[3]) );
	exnor2_3 U223 ( .x(SUM[26]), .a(n61), .b(n98) );
	ao21_3 U224 ( .x(n61), .a(n203), .b(n347), .c(n91) );
	inv_0 U225 ( .x(n62), .a(n166) );
	inv_2 U226 ( .x(n63), .a(n62) );
	nand2_4 U227 ( .x(n166), .a(B[16]), .b(A[16]) );
	inv_0 U228 ( .x(n64), .a(n248) );
	inv_6 U229 ( .x(n248), .a(A[17]) );
	nor2i_2 U23 ( .x(n293), .a(n127), .b(n294) );
	nor2_3 U230 ( .x(n65), .a(A[10]), .b(B[10]) );
	aoai211_1 U231 ( .x(n311), .a(A[0]), .b(n58), .c(n84), .d(n312) );
	nand2i_1 U232 ( .x(n338), .a(A[16]), .b(n247) );
	inv_0 U233 ( .x(n167), .a(n338) );
	inv_0 U234 ( .x(n249), .a(A[18]) );
	nand2_2 U235 ( .x(n133), .a(A[4]), .b(B[4]) );
	exnor2_1 U236 ( .x(SUM[25]), .a(n203), .b(n204) );
	inv_2 U237 ( .x(n68), .a(n293) );
	nand2_0 U238 ( .x(n71), .a(B[9]), .b(A[9]) );
	ao211_5 U239 ( .x(n345), .a(n188), .b(n72), .c(n263), .d(n265) );
	nand2_0 U24 ( .x(n125), .a(A[7]), .b(B[7]) );
	inv_0 U240 ( .x(n72), .a(n189) );
	inv_2 U241 ( .x(n188), .a(A[8]) );
	inv_8 U242 ( .x(n226), .a(A[6]) );
	nand4_3 U243 ( .x(n343), .a(n304), .b(n342), .c(n345), .d(n344) );
	oaoi211_2 U245 ( .x(n80), .a(n83), .b(n82), .c(n343), .d(n81) );
	nor2i_0 U246 ( .x(n288), .a(B[17]), .b(n279) );
	nor2i_3 U247 ( .x(n307), .a(n145), .b(n147) );
	oaoi211_3 U248 ( .x(n74), .a(n80), .b(n78), .c(n77), .d(n75) );
	inv_0 U249 ( .x(n350), .a(n74) );
	inv_1 U25 ( .x(n123), .a(n127) );
	inv_2 U250 ( .x(n75), .a(n336) );
	nand2_2 U251 ( .x(n336), .a(n76), .b(n275) );
	inv_0 U252 ( .x(n76), .a(B[27]) );
	nor2i_3 U253 ( .x(n78), .a(n324), .b(n79) );
	inv_2 U254 ( .x(n81), .a(n357) );
	inv_2 U255 ( .x(n82), .a(n244) );
	inv_2 U256 ( .x(n83), .a(n243) );
	inv_0 U257 ( .x(n275), .a(A[27]) );
	nand2i_2 U258 ( .x(n274), .a(n237), .b(n241) );
	nand2_0 U259 ( .x(n152), .a(A[26]), .b(B[26]) );
	nand2i_2 U26 ( .x(n292), .a(n149), .b(n220) );
	nand2_0 U260 ( .x(n242), .a(B[24]), .b(A[24]) );
	nand2i_2 U261 ( .x(n239), .a(n240), .b(n241) );
	nand2_1 U262 ( .x(n324), .a(n360), .b(A[24]) );
	nand2_0 U264 ( .x(n357), .a(B[23]), .b(A[23]) );
	inv_0 U265 ( .x(n244), .a(B[23]) );
	inv_0 U266 ( .x(n243), .a(A[23]) );
	inv_0 U267 ( .x(n330), .a(n84) );
	inv_2 U268 ( .x(n88), .a(B[7]) );
	nand2i_2 U27 ( .x(n291), .a(n128), .b(n221) );
	inv_0 U270 ( .x(n227), .a(A[7]) );
	inv_0 U271 ( .x(n233), .a(n223) );
	inv_2 U272 ( .x(n91), .a(n237) );
	nand2_0 U273 ( .x(n237), .a(A[25]), .b(B[25]) );
	inv_2 U274 ( .x(n240), .a(n347) );
	exnor2_1 U275 ( .x(n284), .a(B[29]), .b(A[29]) );
	exor2_1 U276 ( .x(n208), .a(A[20]), .b(B[20]) );
	nor2_0 U277 ( .x(n136), .a(A[20]), .b(B[20]) );
	nor2i_3 U278 ( .x(n309), .a(n145), .b(n147) );
	oai21_3 U279 ( .x(n250), .a(A[18]), .b(n164), .c(B[18]) );
	nor2i_1 U28 ( .x(n224), .a(n290), .b(n222) );
	aoi21_1 U280 ( .x(n162), .a(n163), .b(n139), .c(n164) );
	nor2i_0 U281 ( .x(n117), .a(n71), .b(n119) );
	oai21_1 U282 ( .x(n218), .a(n333), .b(n119), .c(n71) );
	nor2i_1 U283 ( .x(n177), .a(n178), .b(n179) );
	inv_0 U284 ( .x(n281), .a(n94) );
	exor2_1 U285 ( .x(SUM[24]), .a(n108), .b(n205) );
	ao21_3 U286 ( .x(n203), .a(n346), .b(n108), .c(n358) );
	aoi21_1 U287 ( .x(n137), .a(n138), .b(n139), .c(n140) );
	ao21_1 U288 ( .x(n193), .a(A[8]), .b(B[8]), .c(n317) );
	nor2_0 U289 ( .x(n187), .a(B[8]), .b(A[8]) );
	or3i_2 U29 ( .x(n222), .a(n223), .b(n219), .c(n114) );
	nand2i_2 U290 ( .x(n264), .a(B[22]), .b(n245) );
	nand2i_3 U291 ( .x(n185), .a(B[11]), .b(n254) );
	inv_2 U292 ( .x(n97), .a(n102) );
	exor2_1 U293 ( .x(SUM[28]), .a(n199), .b(n200) );
	nor2_0 U294 ( .x(n111), .a(A[0]), .b(B[0]) );
	and3i_1 U295 ( .x(n361), .a(n362), .b(B[0]), .c(A[0]) );
	nand2_0 U296 ( .x(n110), .a(A[0]), .b(B[0]) );
	mux2i_1 U297 ( .x(n112), .d0(n288), .sl(n64), .d1(n285) );
	exor2_1 U298 ( .x(n211), .a(B[18]), .b(A[18]) );
	inv_2 U299 ( .x(n98), .a(n151) );
	inv_2 U30 ( .x(n360), .a(n239) );
	nor2i_1 U300 ( .x(n151), .a(n152), .b(n153) );
	inv_0 U301 ( .x(n99), .a(n277) );
	oai21_5 U302 ( .x(n161), .a(n92), .b(n249), .c(n250) );
	nand2_5 U303 ( .x(n344), .a(n143), .b(n264) );
	nor2i_3 U304 ( .x(n100), .a(n337), .b(n261) );
	inv_0 U305 ( .x(n262), .a(n100) );
	inv_0 U306 ( .x(n138), .a(n261) );
	inv_0 U307 ( .x(n101), .a(n343) );
	ao221_4 U308 ( .x(n196), .a(n308), .b(n307), .c(n310), .d(n309), .e(n182) );
	nor2i_3 U309 ( .x(n310), .a(B[30]), .b(n146) );
	inv_2 U31 ( .x(n183), .a(A[30]) );
	and3i_1 U310 ( .x(n144), .a(n147), .b(n145), .c(n352) );
	exnor2_1 U311 ( .x(SUM[22]), .a(n141), .b(n207) );
	nor2_0 U312 ( .x(n163), .a(n94), .b(n167) );
	nand2i_0 U313 ( .x(n145), .a(B[29]), .b(n320) );
	exnor2_3 U314 ( .x(SUM[30]), .a(n144), .b(n282) );
	aoi22_2 U315 ( .x(n304), .a(n299), .b(n305), .c(n306), .d(n303) );
	nor2i_0 U316 ( .x(n141), .a(n142), .b(n143) );
	exnor2_5 U317 ( .x(SUM[31]), .a(n196), .b(n107) );
	inv_2 U318 ( .x(n102), .a(n351) );
	nand2i_0 U319 ( .x(n351), .a(B[28]), .b(n319) );
	nor2i_1 U32 ( .x(n182), .a(B[30]), .b(n183) );
	buf_1 U320 ( .x(n103), .a(n50) );
	inv_0 U321 ( .x(n140), .a(n104) );
	nand2_0 U322 ( .x(n276), .a(A[20]), .b(B[20]) );
	inv_0 U323 ( .x(n253), .a(B[20]) );
	nand2i_0 U324 ( .x(n199), .a(n349), .b(n350) );
	inv_2 U325 ( .x(n107), .a(n197) );
	exor2_1 U326 ( .x(n197), .a(B[31]), .b(A[31]) );
	aoi21_1 U327 ( .x(n160), .a(n66), .b(n139), .c(n99) );
	inv_0 U328 ( .x(n283), .a(n96) );
	nand2i_4 U329 ( .x(n352), .a(A[29]), .b(n96) );
	inv_5 U33 ( .x(n147), .a(n321) );
	nand3i_5 U330 ( .x(n265), .a(n52), .b(n185), .c(n266) );
	nand2i_4 U331 ( .x(n271), .a(n272), .b(n266) );
	nand2_2 U332 ( .x(n297), .a(n298), .b(n169) );
	nor2i_5 U333 ( .x(n299), .a(n300), .b(n263) );
	nand2i_4 U334 ( .x(n278), .a(n252), .b(n161) );
	nand2i_4 U335 ( .x(n216), .a(n184), .b(n340) );
	inv_5 U336 ( .x(n341), .a(n216) );
	oai21_4 U337 ( .x(n215), .a(n341), .b(n176), .c(n175) );
	oai21_4 U338 ( .x(n212), .a(n170), .b(n354), .c(n169) );
	nand3i_3 U339 ( .x(n305), .a(n297), .b(n359), .c(n356) );
	inv_2 U34 ( .x(n256), .a(n300) );
	inv_5 U340 ( .x(n312), .a(n271) );
	nand2_8 U341 ( .x(n181), .a(B[10]), .b(A[10]) );
	nand2_6 U342 ( .x(n175), .a(B[12]), .b(A[12]) );
	nand2_8 U343 ( .x(n348), .a(A[27]), .b(B[27]) );
	nand2i_6 U345 ( .x(n301), .a(A[9]), .b(n232) );
	inv_6 U347 ( .x(n277), .a(n161) );
	nand2_4 U348 ( .x(n342), .a(A[22]), .b(B[22]) );
	inv_0 U35 ( .x(n268), .a(A[15]) );
	inv_6 U352 ( .x(n266), .a(n255) );
	nor2i_2 U353 ( .x(n296), .a(B[8]), .b(n119) );
	nor2_1 U354 ( .x(n365), .a(n366), .b(n231) );
	inv_0 U355 ( .x(n234), .a(n365) );
	inv_0 U356 ( .x(n366), .a(B[2]) );
	inv_3 U357 ( .x(n231), .a(A[2]) );
	nor2i_3 U358 ( .x(n367), .a(n368), .b(A[14]) );
	inv_4 U359 ( .x(n257), .a(n367) );
	aoi22_1 U36 ( .x(n313), .a(n305), .b(n300), .c(n314), .d(n315) );
	inv_0 U360 ( .x(n368), .a(B[14]) );
	nand2i_4 U361 ( .x(n221), .a(B[5]), .b(n228) );
	nand2_2 U362 ( .x(n130), .a(A[5]), .b(B[5]) );
	nand2_3 U363 ( .x(n169), .a(A[14]), .b(B[14]) );
	nand2_1 U364 ( .x(n298), .a(B[15]), .b(A[15]) );
	nand2i_4 U365 ( .x(n122), .a(B[6]), .b(n226) );
	nand2_2 U366 ( .x(n127), .a(A[6]), .b(B[6]) );
	nand2i_0 U367 ( .x(n241), .a(B[26]), .b(n235) );
	nand2_1 U368 ( .x(n323), .a(n360), .b(B[24]) );
	and2_2 U37 ( .x(n58), .a(n224), .b(n57) );
	inv_2 U38 ( .x(n245), .a(A[22]) );
	inv_2 U39 ( .x(n314), .a(n265) );
	nand2_2 U40 ( .x(n263), .a(n100), .b(n264) );
	oai211_1 U41 ( .x(n189), .a(n65), .b(n118), .c(n178), .d(n181) );
	nand2i_2 U42 ( .x(n306), .a(B[8]), .b(n188) );
	nor2i_0 U43 ( .x(n148), .a(n149), .b(n150) );
	inv_2 U44 ( .x(n219), .a(B[0]) );
	nand2i_2 U45 ( .x(n223), .a(B[2]), .b(n231) );
	nor2i_0 U46 ( .x(n126), .a(n127), .b(n128) );
	inv_5 U48 ( .x(n128), .a(n122) );
	nand2_1 U49 ( .x(n192), .a(n330), .b(n331) );
	inv_0 U5 ( .x(n49), .a(n159) );
	nand3i_1 U50 ( .x(n316), .a(n317), .b(n185), .c(n302) );
	or3i_2 U51 ( .x(n340), .a(n192), .b(n119), .c(n316) );
	inv_2 U52 ( .x(n302), .a(n65) );
	inv_2 U53 ( .x(n186), .a(n315) );
	nor3i_1 U54 ( .x(n184), .a(n185), .b(n186), .c(n52) );
	inv_2 U55 ( .x(n294), .a(n125) );
	oai21_1 U56 ( .x(n121), .a(n131), .b(n335), .c(n130) );
	inv_2 U57 ( .x(n131), .a(n221) );
	nand2_2 U58 ( .x(n202), .a(n336), .b(n348) );
	nand2_2 U59 ( .x(n322), .a(n323), .b(n324) );
	inv_2 U6 ( .x(n50), .a(n49) );
	nor2i_1 U60 ( .x(SUM[0]), .a(n110), .b(n111) );
	inv_2 U61 ( .x(n254), .a(A[11]) );
	inv_2 U62 ( .x(n179), .a(n185) );
	nand2_2 U63 ( .x(n178), .a(A[11]), .b(B[11]) );
	oai21_1 U64 ( .x(n217), .a(n65), .b(n355), .c(n181) );
	inv_0 U65 ( .x(n251), .a(A[19]) );
	nand2i_2 U66 ( .x(n260), .a(n135), .b(n66) );
	inv_0 U67 ( .x(n270), .a(B[13]) );
	nand2i_2 U68 ( .x(n258), .a(A[12]), .b(n269) );
	inv_0 U69 ( .x(n269), .a(B[12]) );
	aoai211_3 U7 ( .x(n159), .a(n277), .b(n252), .c(n251), .d(n278) );
	inv_2 U70 ( .x(n339), .a(n175) );
	nor2i_1 U71 ( .x(n180), .a(n181), .b(n65) );
	inv_2 U72 ( .x(n355), .a(n218) );
	exor2_1 U73 ( .x(n207), .a(A[22]), .b(B[22]) );
	nand2i_1 U74 ( .x(n142), .a(n262), .b(n139) );
	exor2_1 U76 ( .x(n210), .a(A[19]), .b(B[19]) );
	oa211_3 U77 ( .x(n66), .a(A[18]), .b(B[18]), .c(n93), .d(n338) );
	inv_0 U78 ( .x(n134), .a(n220) );
	inv_2 U79 ( .x(n229), .a(A[4]) );
	oaoi211_2 U8 ( .x(n104), .a(A[20]), .b(n106), .c(n159), .d(n105) );
	nand2i_2 U80 ( .x(n220), .a(B[4]), .b(n229) );
	nand2i_2 U81 ( .x(n198), .a(n56), .b(n327) );
	nand2i_2 U82 ( .x(n327), .a(n225), .b(n328) );
	inv_0 U83 ( .x(n328), .a(n222) );
	nand2i_2 U84 ( .x(n326), .a(B[3]), .b(n230) );
	inv_0 U85 ( .x(n230), .a(A[3]) );
	nand2i_2 U86 ( .x(n149), .a(n73), .b(B[3]) );
	oai21_2 U87 ( .x(n139), .a(n187), .b(n311), .c(n313) );
	exnor2_1 U88 ( .x(n282), .a(B[30]), .b(A[30]) );
	inv_2 U89 ( .x(n320), .a(A[29]) );
	nor2_0 U9 ( .x(n114), .a(B[1]), .b(A[1]) );
	nand2i_2 U90 ( .x(n325), .a(B[8]), .b(n188) );
	inv_2 U91 ( .x(n67), .a(n295) );
	inv_2 U92 ( .x(n69), .a(n292) );
	inv_2 U93 ( .x(n70), .a(n291) );
	aoi211_1 U94 ( .x(n89), .a(n70), .b(n69), .c(n68), .d(n67) );
	inv_2 U95 ( .x(n85), .a(n56) );
	inv_2 U96 ( .x(n86), .a(n57) );
	oaoi211_1 U97 ( .x(n84), .a(n86), .b(n85), .c(n89), .d(n87) );
	nand2i_2 U98 ( .x(n331), .a(n225), .b(n58) );
	inv_0 U99 ( .x(n225), .a(A[0]) );

endmodule


module EX_DW01_sub_32_0_test_1 (  A, B, CI, DIFF, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] DIFF;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
	n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
	n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
	n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
	n281, n282, n283, n284, n285, n286, n287, n289, n290, n291, n292, n293,
	n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
	n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316, n317,
	n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
	n330, n331, n332, n333, n334, n335, n336, n50, n51, n52, n53, n54, n55,
	n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
	n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
	n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
	n98, n99;


	inv_1 U10 ( .x(n298), .a(n175) );
	exor2_1 U100 ( .x(DIFF[7]), .a(n186), .b(n111) );
	oai21_1 U101 ( .x(n186), .a(n116), .b(n313), .c(n85) );
	inv_2 U102 ( .x(n206), .a(n74) );
	inv_2 U103 ( .x(n313), .a(n187) );
	nor2i_1 U104 ( .x(n111), .a(n112), .b(n113) );
	inv_2 U105 ( .x(n113), .a(n204) );
	exnor2_1 U106 ( .x(DIFF[27]), .a(n194), .b(n195) );
	aoai211_1 U107 ( .x(n194), .a(n329), .b(n328), .c(n272), .d(n327) );
	inv_2 U108 ( .x(n272), .a(n61) );
	inv_2 U109 ( .x(n327), .a(n249) );
	nand2_2 U11 ( .x(n285), .a(n282), .b(n283) );
	nand2_2 U110 ( .x(n195), .a(n314), .b(n130) );
	nand2_2 U111 ( .x(DIFF[0]), .a(n178), .b(n179) );
	inv_2 U112 ( .x(n242), .a(n81) );
	exor2_1 U113 ( .x(DIFF[20]), .a(n332), .b(n147) );
	inv_2 U115 ( .x(n296), .a(n247) );
	nor2_1 U116 ( .x(n147), .a(n126), .b(n148) );
	nor2_1 U117 ( .x(n157), .a(n158), .b(n71) );
	oai21_1 U118 ( .x(n89), .a(n160), .b(n324), .c(n237) );
	exor2_1 U119 ( .x(DIFF[14]), .a(n89), .b(n157) );
	nand2i_2 U12 ( .x(n228), .a(n164), .b(n52) );
	exor2_1 U120 ( .x(DIFF[13]), .a(n201), .b(n159) );
	inv_2 U121 ( .x(n164), .a(n284) );
	nor2_1 U122 ( .x(n159), .a(n160), .b(n161) );
	inv_2 U123 ( .x(n160), .a(n227) );
	inv_2 U124 ( .x(n161), .a(n237) );
	inv_2 U125 ( .x(n324), .a(n201) );
	inv_0 U126 ( .x(n166), .a(n84) );
	nor2_0 U127 ( .x(n165), .a(n81), .b(n166) );
	inv_2 U13 ( .x(n79), .a(n286) );
	exnor2_1 U130 ( .x(DIFF[22]), .a(n127), .b(n141) );
	aoi21_1 U131 ( .x(n127), .a(n51), .b(n125), .c(n128) );
	nor2i_1 U132 ( .x(n141), .a(n142), .b(n143) );
	inv_2 U133 ( .x(n143), .a(n244) );
	exor2_1 U134 ( .x(DIFF[5]), .a(n188), .b(n117) );
	oai21_1 U135 ( .x(n188), .a(n211), .b(n311), .c(n304) );
	inv_2 U136 ( .x(n211), .a(n303) );
	inv_5 U137 ( .x(n311), .a(n189) );
	nor2_1 U138 ( .x(n117), .a(n104), .b(n118) );
	inv_2 U139 ( .x(n104), .a(n305) );
	inv_2 U14 ( .x(n156), .a(n224) );
	inv_2 U140 ( .x(n118), .a(n205) );
	mux2i_1 U141 ( .x(DIFF[19]), .d0(n149), .sl(n91), .d1(n274) );
	aoi21_1 U142 ( .x(n149), .a(A[19]), .b(n150), .c(n151) );
	inv_0 U143 ( .x(n150), .a(B[19]) );
	inv_2 U144 ( .x(n151), .a(n246) );
	exor2_1 U145 ( .x(n274), .a(B[19]), .b(A[19]) );
	exnor2_1 U146 ( .x(DIFF[4]), .a(n189), .b(n190) );
	nand2i_4 U147 ( .x(n189), .a(n180), .b(n309) );
	nand2_2 U148 ( .x(n190), .a(n304), .b(n303) );
	exnor2_1 U149 ( .x(DIFF[18]), .a(n100), .b(n152) );
	oai22_1 U15 ( .x(n291), .a(n223), .b(n237), .c(n156), .d(n236) );
	inv_0 U150 ( .x(n101), .a(n256) );
	nor2_1 U151 ( .x(n152), .a(n153), .b(n94) );
	inv_2 U152 ( .x(n94), .a(n260) );
	nor2i_0 U153 ( .x(n129), .a(n130), .b(n131) );
	exnor2_1 U154 ( .x(n269), .a(A[28]), .b(B[28]) );
	exnor2_1 U155 ( .x(DIFF[8]), .a(n185), .b(n108) );
	inv_2 U156 ( .x(n307), .a(n121) );
	nor2_1 U157 ( .x(n108), .a(n109), .b(n110) );
	inv_2 U158 ( .x(n110), .a(n240) );
	exor2_1 U159 ( .x(n193), .a(B[29]), .b(n58) );
	exor2_1 U160 ( .x(DIFF[29]), .a(n192), .b(n193) );
	exor2_1 U161 ( .x(DIFF[9]), .a(n184), .b(n105) );
	inv_2 U162 ( .x(n109), .a(n231) );
	nor2_1 U163 ( .x(n105), .a(n106), .b(n107) );
	inv_2 U164 ( .x(n106), .a(n239) );
	inv_2 U165 ( .x(n107), .a(n230) );
	inv_2 U166 ( .x(n312), .a(n184) );
	nor2i_1 U167 ( .x(n154), .a(n155), .b(n156) );
	exnor2_1 U168 ( .x(DIFF[17]), .a(n96), .b(n275) );
	inv_2 U169 ( .x(n126), .a(n221) );
	nor2i_1 U170 ( .x(n144), .a(n145), .b(n146) );
	exnor2_1 U171 ( .x(DIFF[23]), .a(n272), .b(n273) );
	exor2_1 U172 ( .x(DIFF[24]), .a(n270), .b(n271) );
	inv_2 U173 ( .x(n215), .a(A[23]) );
	inv_2 U174 ( .x(n140), .a(n216) );
	nor2i_1 U175 ( .x(n138), .a(n139), .b(n140) );
	inv_2 U176 ( .x(n316), .a(n214) );
	inv_2 U177 ( .x(n136), .a(n219) );
	inv_2 U178 ( .x(n137), .a(n251) );
	exor2_1 U179 ( .x(DIFF[3]), .a(n191), .b(n132) );
	inv_2 U180 ( .x(n236), .a(n71) );
	and2_1 U181 ( .x(n50), .a(n216), .b(n217) );
	and3_5 U183 ( .x(n54), .a(n204), .b(n205), .c(n206) );
	ao221_1 U184 ( .x(n56), .a(n296), .b(n53), .c(n128), .d(n244), .e(n297) );
	inv_2 U186 ( .x(n57), .a(n254) );
	inv_2 U187 ( .x(n254), .a(A[30]) );
	inv_2 U188 ( .x(n58), .a(n212) );
	inv_10 U189 ( .x(n131), .a(n317) );
	inv_2 U19 ( .x(n84), .a(n60) );
	nand2i_1 U190 ( .x(n133), .a(B[3]), .b(A[3]) );
	nand2i_2 U191 ( .x(n281), .a(A[3]), .b(B[3]) );
	nand3_1 U192 ( .x(n93), .a(n259), .b(n261), .c(n262) );
	nand2i_6 U193 ( .x(n259), .a(B[17]), .b(n99) );
	nand2i_3 U194 ( .x(n303), .a(A[4]), .b(B[4]) );
	aoi211_1 U195 ( .x(n91), .a(n92), .b(n93), .c(n94), .d(n95) );
	inv_2 U196 ( .x(n153), .a(n92) );
	and3i_1 U197 ( .x(n95), .a(n122), .b(n92), .c(n101) );
	nand2_2 U198 ( .x(n170), .a(n92), .b(n246) );
	nand2_2 U199 ( .x(n245), .a(n92), .b(n246) );
	nand4i_1 U20 ( .x(n229), .a(n119), .b(n84), .c(n230), .d(n231) );
	inv_0 U200 ( .x(n243), .a(A[11]) );
	exnor2_1 U201 ( .x(n277), .a(A[11]), .b(B[11]) );
	nand2i_2 U202 ( .x(n240), .a(B[8]), .b(A[8]) );
	nand2i_2 U203 ( .x(n204), .a(A[7]), .b(B[7]) );
	exnor2_1 U204 ( .x(DIFF[28]), .a(n129), .b(n269) );
	or3i_1 U205 ( .x(n286), .a(n227), .b(n225), .c(n223) );
	inv_2 U208 ( .x(n290), .a(n155) );
	nor2i_2 U209 ( .x(n60), .a(n82), .b(n59) );
	nand2i_2 U21 ( .x(n328), .a(n215), .b(n326) );
	inv_0 U210 ( .x(n59), .a(B[10]) );
	inv_2 U211 ( .x(n82), .a(A[10]) );
	ao211_1 U212 ( .x(n61), .a(n77), .b(n62), .c(n56), .d(n55) );
	nand4_3 U213 ( .x(n62), .a(n287), .b(n292), .c(n73), .d(n330) );
	nand4_1 U214 ( .x(n97), .a(n73), .b(n292), .c(n333), .d(n330) );
	inv_2 U215 ( .x(n122), .a(n97) );
	nand2_1 U216 ( .x(n260), .a(n63), .b(A[18]) );
	inv_0 U217 ( .x(n63), .a(B[18]) );
	nand2i_3 U218 ( .x(n90), .a(A[14]), .b(B[14]) );
	nor2i_1 U219 ( .x(n64), .a(n65), .b(n212) );
	nand2i_2 U22 ( .x(n329), .a(B[23]), .b(n326) );
	inv_0 U220 ( .x(n65), .a(B[29]) );
	nor2_1 U221 ( .x(n66), .a(n212), .b(n67) );
	inv_2 U222 ( .x(n67), .a(n252) );
	ao21_6 U223 ( .x(n68), .a(n182), .b(n183), .c(n131) );
	and2_1 U224 ( .x(n69), .a(n65), .b(n252) );
	ao21_6 U225 ( .x(n70), .a(n182), .b(n183), .c(n131) );
	inv_2 U226 ( .x(n212), .a(A[29]) );
	nand2i_0 U227 ( .x(n252), .a(A[28]), .b(B[28]) );
	nand2i_2 U228 ( .x(n261), .a(B[17]), .b(A[17]) );
	nor3i_2 U229 ( .x(n174), .a(A[17]), .b(B[17]), .c(n175) );
	inv_2 U23 ( .x(n326), .a(n218) );
	nor2i_3 U230 ( .x(n71), .a(n72), .b(n76) );
	inv_0 U231 ( .x(n72), .a(B[14]) );
	aoi31_3 U232 ( .x(n73), .a(n80), .b(n234), .c(n293), .d(n79) );
	exnor2_1 U233 ( .x(n275), .a(B[17]), .b(A[17]) );
	nand2i_0 U234 ( .x(n257), .a(A[17]), .b(B[17]) );
	nand2i_2 U235 ( .x(n295), .a(A[17]), .b(B[17]) );
	nand2i_2 U236 ( .x(n305), .a(B[5]), .b(A[5]) );
	nand2i_2 U237 ( .x(n205), .a(A[5]), .b(B[5]) );
	nor2_3 U238 ( .x(n74), .a(A[6]), .b(n75) );
	nand2_2 U239 ( .x(n85), .a(n75), .b(A[6]) );
	nand2_2 U24 ( .x(n218), .a(n50), .b(n219) );
	inv_0 U240 ( .x(n158), .a(n90) );
	inv_0 U241 ( .x(n76), .a(A[14]) );
	nand2i_0 U242 ( .x(n179), .a(B[0]), .b(A[0]) );
	nand2i_2 U243 ( .x(n92), .a(A[18]), .b(B[18]) );
	ao211_5 U244 ( .x(n315), .a(n77), .b(n62), .c(n56), .d(n55) );
	nand4i_1 U245 ( .x(n294), .a(n245), .b(n53), .c(n98), .d(n295) );
	exnor2_1 U246 ( .x(n271), .a(A[24]), .b(B[24]) );
	nand2i_2 U247 ( .x(n217), .a(A[24]), .b(B[24]) );
	nand2i_2 U249 ( .x(n320), .a(B[30]), .b(n253) );
	nand2i_2 U25 ( .x(n247), .a(B[19]), .b(A[19]) );
	exnor2_3 U250 ( .x(DIFF[31]), .a(n266), .b(n78) );
	inv_2 U251 ( .x(n78), .a(n267) );
	exnor2_1 U252 ( .x(n267), .a(A[31]), .b(B[31]) );
	nand2i_2 U253 ( .x(n231), .a(A[8]), .b(B[8]) );
	nand2i_3 U254 ( .x(n239), .a(B[9]), .b(A[9]) );
	aoai211_1 U255 ( .x(n172), .a(n182), .b(n183), .c(n131), .d(n69) );
	aoai211_1 U256 ( .x(n173), .a(n182), .b(n183), .c(n131), .d(n66) );
	aoai211_1 U257 ( .x(n192), .a(n182), .b(n183), .c(n131), .d(n252) );
	or2_6 U258 ( .x(n80), .a(n120), .b(n121) );
	inv_4 U259 ( .x(n293), .a(n228) );
	aoi21_1 U26 ( .x(n167), .a(n168), .b(n169), .c(n170) );
	exnor2_1 U260 ( .x(DIFF[16]), .a(n97), .b(n200) );
	aoi21_1 U262 ( .x(n96), .a(n97), .b(n98), .c(n99) );
	aoi21_1 U263 ( .x(n100), .a(n101), .b(n97), .c(n93) );
	inv_0 U264 ( .x(n116), .a(n206) );
	nor2i_3 U265 ( .x(n81), .a(n83), .b(n82) );
	inv_0 U266 ( .x(n83), .a(B[10]) );
	nand2i_4 U267 ( .x(n222), .a(A[21]), .b(B[21]) );
	nand2i_2 U268 ( .x(n98), .a(A[16]), .b(B[16]) );
	nand2i_2 U269 ( .x(n227), .a(A[13]), .b(B[13]) );
	nor2i_1 U27 ( .x(n168), .a(n261), .b(n299) );
	nand2i_3 U271 ( .x(n284), .a(A[12]), .b(B[12]) );
	nand2i_2 U272 ( .x(n225), .a(B[12]), .b(A[12]) );
	nand2_2 U273 ( .x(DIFF[1]), .a(n86), .b(n87) );
	aoi21_3 U274 ( .x(n88), .a(n89), .b(n90), .c(n71) );
	nor2_5 U275 ( .x(n102), .a(n103), .b(n104) );
	nor2i_5 U276 ( .x(n119), .a(B[11]), .b(A[11]) );
	aoi21_3 U277 ( .x(n123), .a(n124), .b(n332), .c(n126) );
	nor2_5 U278 ( .x(n135), .a(n136), .b(n137) );
	and3i_3 U279 ( .x(n171), .a(n64), .b(n172), .c(n173) );
	inv_0 U28 ( .x(n169), .a(n258) );
	exor2_3 U280 ( .x(DIFF[26]), .a(n196), .b(n135) );
	exor2_3 U281 ( .x(DIFF[25]), .a(n197), .b(n138) );
	exnor2_3 U282 ( .x(DIFF[21]), .a(n123), .b(n144) );
	exnor2_5 U283 ( .x(DIFF[15]), .a(n88), .b(n154) );
	aoai211_4 U285 ( .x(n238), .a(n239), .b(n240), .c(n241), .d(n242) );
	aoai211_4 U286 ( .x(n263), .a(n264), .b(B[11]), .c(n243), .d(n265) );
	exnor2_5 U287 ( .x(DIFF[30]), .a(n171), .b(n268) );
	exor2_3 U288 ( .x(DIFF[11]), .a(n276), .b(n277) );
	aoi21_3 U289 ( .x(n292), .a(n293), .b(n263), .c(n291) );
	nand2_2 U29 ( .x(n258), .a(n259), .b(n260) );
	nand2i_4 U290 ( .x(n304), .a(B[4]), .b(A[4]) );
	oai211_4 U291 ( .x(n310), .a(n311), .b(n210), .c(n307), .d(n306) );
	oai21_4 U292 ( .x(n184), .a(n185), .b(n109), .c(n240) );
	nand2i_4 U293 ( .x(n314), .a(A[27]), .b(B[27]) );
	inv_5 U294 ( .x(n264), .a(n238) );
	aoai211_4 U295 ( .x(n317), .a(n318), .b(n315), .c(n249), .d(n314) );
	inv_5 U296 ( .x(n323), .a(n202) );
	oai21_4 U297 ( .x(n201), .a(n164), .b(n323), .c(n225) );
	inv_5 U298 ( .x(n325), .a(n203) );
	oai21_4 U299 ( .x(n276), .a(n166), .b(n325), .c(n242) );
	nand2i_2 U30 ( .x(n244), .a(A[22]), .b(B[22]) );
	aoai211_4 U300 ( .x(n270), .a(B[23]), .b(n215), .c(n272), .d(n220) );
	exnor2_3 U301 ( .x(n268), .a(n57), .b(B[30]) );
	nand2i_5 U302 ( .x(n202), .a(n263), .b(n322) );
	ao21_4 U303 ( .x(n197), .a(n217), .b(n270), .c(n316) );
	ao21_4 U304 ( .x(n196), .a(n50), .b(n270), .c(n255) );
	inv_6 U305 ( .x(n185), .a(n310) );
	nand2i_5 U306 ( .x(n322), .a(n229), .b(n310) );
	or3i_5 U307 ( .x(n330), .a(n334), .b(n285), .c(n279) );
	nand2i_6 U308 ( .x(n282), .a(A[2]), .b(B[2]) );
	nor2i_5 U309 ( .x(n180), .a(n178), .b(n181) );
	nand2i_0 U31 ( .x(n142), .a(B[22]), .b(A[22]) );
	nand2i_4 U310 ( .x(n265), .a(B[11]), .b(n238) );
	nand2i_6 U311 ( .x(n224), .a(A[15]), .b(B[15]) );
	nand2i_8 U312 ( .x(n246), .a(A[19]), .b(B[19]) );
	nand2i_6 U313 ( .x(n210), .a(n211), .b(n54) );
	nand2i_5 U314 ( .x(n306), .a(n102), .b(n54) );
	nand2_6 U315 ( .x(n223), .a(n224), .b(n90) );
	nand2i_6 U316 ( .x(n175), .a(n170), .b(n53) );
	exnor2_1 U317 ( .x(DIFF[10]), .a(n203), .b(n331) );
	inv_2 U318 ( .x(n331), .a(n165) );
	oai21_2 U319 ( .x(n203), .a(n312), .b(n107), .c(n239) );
	oai21_1 U32 ( .x(n128), .a(n146), .b(n221), .c(n145) );
	or3i_3 U320 ( .x(n332), .a(n300), .b(n296), .c(n167) );
	or3i_3 U321 ( .x(n300), .a(n97), .b(n245), .c(n256) );
	or3i_1 U322 ( .x(n125), .a(n300), .b(n296), .c(n167) );
	and4_5 U323 ( .x(n334), .a(n335), .b(n234), .c(n52), .d(n235) );
	buf_1 U324 ( .x(n333), .a(n287) );
	aoi21_3 U325 ( .x(n287), .a(n334), .b(n336), .c(n290) );
	inv_2 U326 ( .x(n335), .a(n233) );
	inv_6 U327 ( .x(n234), .a(n229) );
	inv_4 U328 ( .x(n235), .a(n210) );
	and2_5 U329 ( .x(n52), .a(n226), .b(n227) );
	inv_0 U33 ( .x(n146), .a(n222) );
	nand2_0 U330 ( .x(n233), .a(n284), .b(n281) );
	and2_6 U331 ( .x(n53), .a(n51), .b(n244) );
	and2_5 U332 ( .x(n51), .a(n124), .b(n222) );
	aoai211_2 U333 ( .x(n266), .a(B[30]), .b(n319), .c(n254), .d(n320) );
	inv_5 U334 ( .x(n319), .a(n253) );
	oai211_1 U335 ( .x(n336), .a(n308), .b(n208), .c(n133), .d(n301) );
	oai211_1 U336 ( .x(n289), .a(n308), .b(n208), .c(n133), .d(n301) );
	nand2i_0 U337 ( .x(n237), .a(B[13]), .b(A[13]) );
	nand2i_0 U34 ( .x(n221), .a(B[20]), .b(A[20]) );
	inv_0 U35 ( .x(n148), .a(n124) );
	nand2i_2 U36 ( .x(n124), .a(A[20]), .b(B[20]) );
	nand2i_2 U38 ( .x(n309), .a(n134), .b(n289) );
	nand3_1 U39 ( .x(n181), .a(n281), .b(n282), .c(n283) );
	inv_4 U4 ( .x(n226), .a(n223) );
	nand2i_5 U40 ( .x(n178), .a(A[0]), .b(B[0]) );
	nand2_2 U41 ( .x(n256), .a(n98), .b(n257) );
	inv_2 U42 ( .x(n299), .a(n262) );
	inv_2 U43 ( .x(n177), .a(A[17]) );
	nand2i_2 U44 ( .x(n262), .a(n177), .b(n99) );
	oai21_1 U45 ( .x(n121), .a(n113), .b(n85), .c(n112) );
	inv_2 U46 ( .x(n75), .a(B[6]) );
	nand2i_0 U47 ( .x(n112), .a(B[7]), .b(A[7]) );
	inv_2 U48 ( .x(n103), .a(n304) );
	inv_4 U49 ( .x(n120), .a(n306) );
	oai211_1 U51 ( .x(n249), .a(n218), .b(n220), .c(n250), .d(n251) );
	nand2_2 U52 ( .x(n318), .a(n329), .b(n328) );
	nand2i_2 U53 ( .x(n183), .a(n213), .b(n130) );
	inv_2 U54 ( .x(n213), .a(B[28]) );
	nand2i_0 U55 ( .x(n130), .a(B[27]), .b(A[27]) );
	nand2i_2 U56 ( .x(n182), .a(A[28]), .b(n130) );
	ao221_4 U57 ( .x(n253), .a(n70), .b(n69), .c(n68), .d(n66), .e(n64) );
	inv_2 U58 ( .x(n279), .a(n178) );
	nand2i_2 U59 ( .x(n208), .a(B[1]), .b(A[1]) );
	nand2_2 U6 ( .x(n241), .a(n84), .b(n230) );
	inv_2 U60 ( .x(n302), .a(n208) );
	nand2_2 U61 ( .x(n87), .a(n302), .b(n178) );
	nor2i_1 U62 ( .x(n280), .a(B[1]), .b(n178) );
	inv_2 U63 ( .x(n209), .a(B[1]) );
	exnor2_1 U64 ( .x(n278), .a(n279), .b(n209) );
	mux2i_1 U65 ( .x(n86), .d0(n278), .sl(A[1]), .d1(n280) );
	nand2i_2 U66 ( .x(n230), .a(A[9]), .b(B[9]) );
	nand2i_0 U67 ( .x(n155), .a(B[15]), .b(A[15]) );
	nand2i_2 U68 ( .x(n248), .a(B[16]), .b(A[16]) );
	nand2_0 U69 ( .x(n200), .a(n248), .b(n98) );
	nand2i_2 U7 ( .x(n283), .a(A[1]), .b(B[1]) );
	inv_2 U70 ( .x(n99), .a(n248) );
	nand2i_0 U71 ( .x(n145), .a(B[21]), .b(A[21]) );
	exnor2_1 U72 ( .x(n273), .a(A[23]), .b(B[23]) );
	inv_2 U73 ( .x(n77), .a(n294) );
	inv_2 U74 ( .x(n297), .a(n142) );
	ao211_2 U75 ( .x(n55), .a(n298), .b(n258), .c(n174), .d(n176) );
	nand2i_2 U76 ( .x(n220), .a(B[23]), .b(A[23]) );
	nand2i_2 U77 ( .x(n251), .a(B[26]), .b(A[26]) );
	nand2i_2 U78 ( .x(n219), .a(A[26]), .b(B[26]) );
	oai21_1 U79 ( .x(n255), .a(n140), .b(n214), .c(n139) );
	nand2_2 U8 ( .x(n250), .a(n255), .b(n219) );
	nand2i_0 U80 ( .x(n214), .a(B[24]), .b(A[24]) );
	nand2i_2 U81 ( .x(n139), .a(B[25]), .b(A[25]) );
	nand2i_2 U82 ( .x(n216), .a(A[25]), .b(B[25]) );
	inv_2 U83 ( .x(n134), .a(n281) );
	nor2i_1 U84 ( .x(n132), .a(n133), .b(n134) );
	nand2i_2 U85 ( .x(n301), .a(B[2]), .b(A[2]) );
	inv_2 U86 ( .x(n308), .a(n282) );
	oai21_1 U87 ( .x(n191), .a(n308), .b(n321), .c(n301) );
	inv_2 U88 ( .x(n321), .a(n198) );
	nand2_2 U89 ( .x(n199), .a(n282), .b(n301) );
	nor3i_1 U9 ( .x(n176), .a(n99), .b(n177), .c(n175) );
	inv_2 U90 ( .x(n207), .a(A[1]) );
	aoai211_1 U91 ( .x(n198), .a(B[1]), .b(n207), .c(n279), .d(n208) );
	exnor2_1 U92 ( .x(DIFF[2]), .a(n198), .b(n199) );
	exor2_1 U93 ( .x(DIFF[6]), .a(n187), .b(n114) );
	ao21_1 U94 ( .x(n187), .a(n188), .b(n205), .c(n104) );
	nor2_1 U95 ( .x(n114), .a(n115), .b(n116) );
	inv_2 U96 ( .x(n115), .a(n85) );
	exor2_1 U97 ( .x(DIFF[12]), .a(n202), .b(n162) );
	nor2_1 U98 ( .x(n162), .a(n163), .b(n164) );
	inv_2 U99 ( .x(n163), .a(n225) );

endmodule


module EX_DW01_sub_32_1_test_1 (  A, B, CI, DIFF, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] DIFF;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
	n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
	n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
	n280, n281, n282, n283, n284, n50, n51, n52, n53, n54, n55, n56, n57,
	n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71,
	n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
	n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	inv_4 U10 ( .x(n102), .a(n258) );
	nand2i_2 U100 ( .x(n282), .a(n254), .b(n230) );
	and3i_1 U101 ( .x(n151), .a(n154), .b(n152), .c(n52) );
	nand3i_1 U102 ( .x(n166), .a(n151), .b(n258), .c(n282) );
	inv_2 U103 ( .x(n82), .a(n88) );
	inv_0 U104 ( .x(n87), .a(A[22]) );
	aoai211_1 U105 ( .x(DIFF[22]), .a(n85), .b(n86), .c(n87), .d(n88) );
	inv_2 U106 ( .x(n118), .a(n174) );
	inv_2 U107 ( .x(n117), .a(n179) );
	nor2_1 U108 ( .x(n116), .a(n117), .b(n118) );
	ao21_1 U109 ( .x(n159), .a(n269), .b(n160), .c(n121) );
	nand2_2 U11 ( .x(n187), .a(n188), .b(n189) );
	nand2i_2 U110 ( .x(n269), .a(A[4]), .b(B[4]) );
	inv_2 U111 ( .x(n272), .a(n159) );
	nand2i_0 U112 ( .x(n96), .a(n182), .b(n91) );
	inv_0 U113 ( .x(n95), .a(A[19]) );
	aoai211_1 U114 ( .x(DIFF[19]), .a(n93), .b(n94), .c(n95), .d(n96) );
	nor2_1 U115 ( .x(n119), .a(n120), .b(n121) );
	inv_2 U116 ( .x(n121), .a(n262) );
	nand2i_0 U117 ( .x(n262), .a(B[4]), .b(A[4]) );
	inv_2 U118 ( .x(n266), .a(n205) );
	aoai211_1 U119 ( .x(n267), .a(n260), .b(n268), .c(n171), .d(n207) );
	nand2i_2 U12 ( .x(n202), .a(n130), .b(n178) );
	nand4i_1 U120 ( .x(n205), .a(n100), .b(n69), .c(n206), .d(n207) );
	nand2i_3 U121 ( .x(n75), .a(n215), .b(n91) );
	nand2i_2 U122 ( .x(n79), .a(n246), .b(n91) );
	oai211_1 U123 ( .x(DIFF[28]), .a(n73), .b(n74), .c(n75), .d(n76) );
	exor2_1 U124 ( .x(DIFF[8]), .a(n158), .b(n104) );
	nand2_2 U125 ( .x(n158), .a(n155), .b(n270) );
	nor2_0 U126 ( .x(n104), .a(n105), .b(n106) );
	nand2i_3 U127 ( .x(n72), .a(n216), .b(A[29]) );
	nand2_1 U128 ( .x(DIFF[29]), .a(n71), .b(n72) );
	inv_2 U129 ( .x(n128), .a(A[30]) );
	nand2i_2 U13 ( .x(n263), .a(n150), .b(n260) );
	oai21_1 U130 ( .x(DIFF[1]), .a(A[1]), .b(n67), .c(n68) );
	exnor2_1 U131 ( .x(n67), .a(n69), .b(n168) );
	inv_2 U132 ( .x(n168), .a(B[1]) );
	mux2i_1 U133 ( .x(n68), .d0(n260), .sl(n265), .d1(n238) );
	inv_2 U134 ( .x(n260), .a(n170) );
	inv_2 U135 ( .x(n265), .a(n69) );
	nor2_0 U136 ( .x(n101), .a(n102), .b(n103) );
	inv_2 U137 ( .x(n279), .a(n271) );
	inv_2 U138 ( .x(n105), .a(n231) );
	inv_2 U139 ( .x(n152), .a(n176) );
	nor2i_0 U14 ( .x(n150), .a(B[2]), .b(A[2]) );
	nand2_2 U140 ( .x(n255), .a(n55), .b(B[8]) );
	inv_5 U141 ( .x(n106), .a(n255) );
	oai211_1 U142 ( .x(n157), .a(n106), .b(n155), .c(n231), .d(n271) );
	inv_2 U143 ( .x(n199), .a(n259) );
	inv_2 U144 ( .x(n141), .a(n186) );
	inv_2 U145 ( .x(n126), .a(n275) );
	inv_2 U146 ( .x(n125), .a(n224) );
	aoi21_1 U147 ( .x(n252), .a(n125), .b(n189), .c(n126) );
	nand2_2 U148 ( .x(n251), .a(n188), .b(n189) );
	oai21_1 U149 ( .x(n277), .a(n139), .b(n137), .c(n140) );
	nor3_0 U15 ( .x(n185), .a(A[22]), .b(A[20]), .c(A[21]) );
	aoai211_1 U150 ( .x(n163), .a(n186), .b(n277), .c(n251), .d(n252) );
	exor2_1 U151 ( .x(DIFF[16]), .a(n235), .b(n98) );
	inv_2 U152 ( .x(n93), .a(n97) );
	inv_0 U153 ( .x(n122), .a(A[17]) );
	nor2i_1 U154 ( .x(n99), .a(n122), .b(n93) );
	inv_0 U155 ( .x(n98), .a(A[16]) );
	nand4_1 U156 ( .x(n97), .a(n222), .b(n219), .c(n220), .d(n223) );
	aoi31_1 U157 ( .x(DIFF[17]), .a(n97), .b(n98), .c(n91), .d(n99) );
	nand4i_1 U158 ( .x(n90), .a(A[20]), .b(n219), .c(n220), .d(n221) );
	inv_2 U159 ( .x(n83), .a(A[23]) );
	nor2_1 U16 ( .x(n243), .a(A[25]), .b(A[24]) );
	nand4_2 U160 ( .x(n208), .a(n60), .b(n209), .c(n210), .d(n211) );
	nand2i_2 U161 ( .x(n248), .a(A[23]), .b(n214) );
	nand2_2 U162 ( .x(DIFF[25]), .a(n80), .b(n81) );
	oai21_1 U163 ( .x(n81), .a(n53), .b(n247), .c(A[25]) );
	inv_2 U164 ( .x(n78), .a(A[26]) );
	inv_2 U165 ( .x(n77), .a(n80) );
	oai21_1 U166 ( .x(DIFF[26]), .a(n77), .b(n78), .c(n79) );
	exor2_1 U167 ( .x(DIFF[2]), .a(n162), .b(n132) );
	exor2_1 U168 ( .x(DIFF[6]), .a(n108), .b(n114) );
	exnor2_1 U169 ( .x(DIFF[12]), .a(n135), .b(n146) );
	inv_4 U17 ( .x(n56), .a(A[9]) );
	exnor2_1 U170 ( .x(DIFF[7]), .a(n107), .b(n111) );
	exnor2_1 U171 ( .x(DIFF[27]), .a(n73), .b(n218) );
	inv_2 U172 ( .x(n73), .a(n79) );
	inv_0 U173 ( .x(n218), .a(A[27]) );
	exor2_1 U174 ( .x(DIFF[11]), .a(n236), .b(n237) );
	inv_1 U175 ( .x(n89), .a(n182) );
	aoi31_1 U176 ( .x(DIFF[20]), .a(n89), .b(n90), .c(n91), .d(n92) );
	exor2_1 U177 ( .x(DIFF[14]), .a(n165), .b(n142) );
	exnor2_1 U178 ( .x(DIFF[13]), .a(n138), .b(n144) );
	exnor2_1 U179 ( .x(DIFF[10]), .a(n166), .b(n167) );
	nor2_0 U18 ( .x(n253), .a(n106), .b(n103) );
	exor2_1 U180 ( .x(DIFF[5]), .a(n159), .b(n116) );
	exor2_1 U181 ( .x(DIFF[4]), .a(n160), .b(n119) );
	inv_2 U182 ( .x(n94), .a(A[18]) );
	exnor2_1 U183 ( .x(DIFF[18]), .a(n93), .b(n94) );
	exor2_1 U184 ( .x(DIFF[9]), .a(n157), .b(n101) );
	exnor2_1 U185 ( .x(DIFF[15]), .a(n163), .b(n164) );
	inv_2 U186 ( .x(n86), .a(A[21]) );
	exnor2_1 U187 ( .x(DIFF[21]), .a(n85), .b(n86) );
	exnor2_1 U188 ( .x(DIFF[24]), .a(n233), .b(n234) );
	inv_2 U189 ( .x(n233), .a(n84) );
	nand2_3 U19 ( .x(n191), .a(n153), .b(n192) );
	inv_2 U190 ( .x(n234), .a(A[24]) );
	inv_2 U191 ( .x(n232), .a(A[31]) );
	and2_6 U192 ( .x(n50), .a(n195), .b(n140) );
	nand2i_2 U193 ( .x(n281), .a(A[4]), .b(B[4]) );
	inv_2 U194 ( .x(n120), .a(n269) );
	inv_2 U195 ( .x(n177), .a(n280) );
	and2_1 U196 ( .x(n51), .a(n264), .b(n263) );
	inv_0 U197 ( .x(n74), .a(A[28]) );
	nand2_0 U198 ( .x(n76), .a(A[27]), .b(A[28]) );
	inv_2 U199 ( .x(n217), .a(A[29]) );
	nand2_2 U20 ( .x(n230), .a(n155), .b(n231) );
	nand2_8 U200 ( .x(n71), .a(n216), .b(n217) );
	inv_10 U201 ( .x(n216), .a(n75) );
	nor2_0 U202 ( .x(n183), .a(A[18]), .b(A[19]) );
	inv_2 U203 ( .x(n52), .a(n103) );
	inv_0 U204 ( .x(n103), .a(n153) );
	aoi21_5 U205 ( .x(n155), .a(n181), .b(n175), .c(n148) );
	inv_7 U206 ( .x(n273), .a(n201) );
	nand2i_0 U207 ( .x(n261), .a(B[7]), .b(A[7]) );
	nand2i_2 U208 ( .x(n175), .a(A[7]), .b(B[7]) );
	ao21_6 U209 ( .x(n180), .a(n181), .b(n175), .c(n148) );
	inv_2 U21 ( .x(n55), .a(A[8]) );
	inv_2 U210 ( .x(n53), .a(n91) );
	nand2_2 U211 ( .x(n186), .a(n54), .b(A[12]) );
	inv_0 U212 ( .x(n54), .a(B[12]) );
	nand2_4 U213 ( .x(n153), .a(n56), .b(B[9]) );
	inv_0 U214 ( .x(n57), .a(n109) );
	inv_2 U215 ( .x(n58), .a(n57) );
	nand2i_0 U216 ( .x(n174), .a(A[5]), .b(B[5]) );
	nand2i_4 U217 ( .x(n179), .a(B[5]), .b(A[5]) );
	oai211_4 U218 ( .x(n149), .a(n59), .b(A[5]), .c(n58), .d(n175) );
	inv_4 U219 ( .x(n59), .a(B[5]) );
	nand2_0 U22 ( .x(n254), .a(n52), .b(n255) );
	aoai211_3 U220 ( .x(n211), .a(n50), .b(n225), .c(n241), .d(n259) );
	nand2i_2 U221 ( .x(n69), .a(A[0]), .b(B[0]) );
	nand2i_0 U222 ( .x(n70), .a(B[0]), .b(A[0]) );
	inv_2 U223 ( .x(n193), .a(n61) );
	inv_0 U224 ( .x(n62), .a(B[10]) );
	nand2i_4 U225 ( .x(n172), .a(B[3]), .b(A[3]) );
	aoi21_1 U226 ( .x(n107), .a(n108), .b(n58), .c(n110) );
	inv_2 U227 ( .x(n115), .a(n58) );
	nand2i_3 U228 ( .x(n231), .a(B[8]), .b(A[8]) );
	inv_0 U229 ( .x(n64), .a(B[10]) );
	nand2i_0 U23 ( .x(n154), .a(n106), .b(n160) );
	inv_0 U230 ( .x(n65), .a(A[10]) );
	nand2_0 U231 ( .x(n109), .a(n66), .b(B[6]) );
	nand2i_3 U232 ( .x(n189), .a(A[14]), .b(B[14]) );
	nand2i_2 U233 ( .x(n188), .a(A[13]), .b(B[13]) );
	nand2i_4 U234 ( .x(n140), .a(A[12]), .b(B[12]) );
	nand2i_0 U235 ( .x(n257), .a(B[6]), .b(A[6]) );
	oai21_4 U236 ( .x(DIFF[23]), .a(n82), .b(n83), .c(n84) );
	nor2i_5 U237 ( .x(n127), .a(n128), .b(n71) );
	nor3i_5 U238 ( .x(n148), .a(A[4]), .b(B[4]), .c(n149) );
	nand2_5 U239 ( .x(n196), .a(n197), .b(n198) );
	inv_0 U24 ( .x(n264), .a(n171) );
	nand2i_4 U240 ( .x(n201), .a(n202), .b(n203) );
	nand2i_4 U241 ( .x(n204), .a(n149), .b(n203) );
	oai211_3 U242 ( .x(n225), .a(n191), .b(n226), .c(n227), .d(n228) );
	exnor2_5 U243 ( .x(DIFF[31]), .a(n127), .b(n232) );
	exnor2_3 U244 ( .x(DIFF[30]), .a(A[30]), .b(n71) );
	nand4_1 U246 ( .x(n235), .a(n211), .b(n256), .c(n220), .d(n219) );
	inv_5 U247 ( .x(n198), .a(n191) );
	or3i_5 U248 ( .x(n219), .a(n273), .b(n51), .c(n177) );
	or3i_5 U249 ( .x(n220), .a(n274), .b(n177), .c(n205) );
	nand2i_4 U250 ( .x(n242), .a(B[15]), .b(A[15]) );
	nand2_5 U251 ( .x(n256), .a(n203), .b(n180) );
	nand2i_4 U252 ( .x(n80), .a(n212), .b(n91) );
	nand2i_4 U253 ( .x(n88), .a(n184), .b(n91) );
	nand2i_4 U254 ( .x(n84), .a(n248), .b(n91) );
	nand2_2 U255 ( .x(n164), .a(n242), .b(n259) );
	inv_5 U256 ( .x(n274), .a(n204) );
	nand3_3 U257 ( .x(n209), .a(n274), .b(n281), .c(n266) );
	inv_12 U258 ( .x(n91), .a(n208) );
	nand2_8 U259 ( .x(n160), .a(n205), .b(n267) );
	nand2_2 U26 ( .x(n171), .a(n172), .b(n173) );
	nand2i_5 U260 ( .x(n259), .a(A[15]), .b(B[15]) );
	nor3i_5 U261 ( .x(n221), .a(n89), .b(n249), .c(n250) );
	nand3i_5 U262 ( .x(n271), .a(n106), .b(n160), .c(n152) );
	inv_6 U263 ( .x(n203), .a(n156) );
	nand2i_6 U264 ( .x(n206), .a(A[2]), .b(B[2]) );
	nand2i_4 U265 ( .x(n213), .a(A[23]), .b(n243) );
	oai21_5 U266 ( .x(n226), .a(n102), .b(n105), .c(n240) );
	nand3i_5 U267 ( .x(n156), .a(n199), .b(n50), .c(n200) );
	nand2i_5 U268 ( .x(n192), .a(A[11]), .b(B[11]) );
	and2_2 U269 ( .x(n283), .a(n284), .b(A[2]) );
	nand2i_0 U27 ( .x(n268), .a(A[2]), .b(B[2]) );
	inv_2 U270 ( .x(n173), .a(n283) );
	inv_2 U271 ( .x(n284), .a(B[2]) );
	inv_4 U272 ( .x(n240), .a(n63) );
	nor2_3 U273 ( .x(n197), .a(n106), .b(n63) );
	nor2i_3 U274 ( .x(n63), .a(n65), .b(n64) );
	nand2i_2 U28 ( .x(n207), .a(A[3]), .b(B[3]) );
	nor2i_0 U29 ( .x(n100), .a(B[1]), .b(A[1]) );
	nand2i_2 U30 ( .x(n212), .a(n213), .b(n214) );
	inv_2 U31 ( .x(n245), .a(n212) );
	nor2_0 U32 ( .x(n244), .a(A[26]), .b(A[27]) );
	nand3i_1 U33 ( .x(n215), .a(A[28]), .b(n244), .c(n245) );
	nand2i_0 U34 ( .x(n176), .a(n177), .b(n178) );
	nand2_2 U35 ( .x(n270), .a(n152), .b(n160) );
	nor2i_1 U36 ( .x(n238), .a(B[1]), .b(n169) );
	inv_2 U37 ( .x(n178), .a(n149) );
	nor2_1 U38 ( .x(n239), .a(n110), .b(n113) );
	oai21_3 U39 ( .x(n181), .a(n149), .b(n179), .c(n239) );
	nor2_1 U4 ( .x(n124), .a(n125), .b(n126) );
	nor2_1 U40 ( .x(n223), .a(n250), .b(n249) );
	inv_5 U41 ( .x(n250), .a(n211) );
	nor2_0 U42 ( .x(n222), .a(A[16]), .b(A[17]) );
	inv_2 U43 ( .x(n249), .a(n256) );
	nand2i_2 U44 ( .x(n280), .a(A[4]), .b(B[4]) );
	oai221_1 U45 ( .x(n241), .a(n143), .b(n124), .c(n186), .d(n187), .e(n242) );
	inv_2 U46 ( .x(n195), .a(n187) );
	or3i_3 U47 ( .x(n210), .a(n273), .b(n120), .c(n51) );
	inv_2 U48 ( .x(n200), .a(n196) );
	or2_2 U49 ( .x(n60), .a(n155), .b(n156) );
	nand2i_2 U5 ( .x(n228), .a(n194), .b(n61) );
	nand3i_0 U50 ( .x(n247), .a(A[23]), .b(n234), .c(n214) );
	nand2i_2 U51 ( .x(n184), .a(n182), .b(n185) );
	nand2i_0 U52 ( .x(n246), .a(A[26]), .b(n245) );
	inv_2 U53 ( .x(n214), .a(n184) );
	exor2_1 U54 ( .x(DIFF[3]), .a(n161), .b(n129) );
	oai21_1 U55 ( .x(n161), .a(n134), .b(n276), .c(n133) );
	nor2_1 U56 ( .x(n129), .a(n130), .b(n131) );
	inv_2 U57 ( .x(n130), .a(n207) );
	inv_0 U58 ( .x(n131), .a(n172) );
	inv_2 U59 ( .x(n134), .a(n206) );
	inv_2 U6 ( .x(n194), .a(A[11]) );
	nand2i_0 U60 ( .x(n133), .a(B[2]), .b(A[2]) );
	nor2i_1 U61 ( .x(n132), .a(n133), .b(n134) );
	aoai211_1 U62 ( .x(n162), .a(B[1]), .b(n169), .c(n265), .d(n170) );
	inv_2 U63 ( .x(n169), .a(A[1]) );
	nand2i_2 U64 ( .x(n170), .a(B[1]), .b(A[1]) );
	inv_2 U65 ( .x(n276), .a(n162) );
	nor2_1 U66 ( .x(n114), .a(n110), .b(n115) );
	nor2_1 U67 ( .x(n146), .a(n141), .b(n147) );
	nand4_1 U68 ( .x(n136), .a(n200), .b(n178), .c(n280), .d(n160) );
	nor2i_1 U69 ( .x(n135), .a(n136), .b(n137) );
	nor2i_0 U7 ( .x(n61), .a(n62), .b(n65) );
	nor2_1 U70 ( .x(n111), .a(n112), .b(n113) );
	inv_2 U71 ( .x(n112), .a(n175) );
	inv_2 U72 ( .x(n113), .a(n261) );
	oai21_1 U73 ( .x(n108), .a(n118), .b(n272), .c(n179) );
	inv_0 U74 ( .x(n66), .a(A[6]) );
	inv_2 U75 ( .x(n110), .a(n257) );
	nand2_2 U76 ( .x(DIFF[0]), .a(n69), .b(n70) );
	exnor2_1 U77 ( .x(n237), .a(B[11]), .b(A[11]) );
	oai21_1 U79 ( .x(n278), .a(n279), .b(n230), .c(n253) );
	inv_0 U8 ( .x(n190), .a(B[11]) );
	nand2i_2 U80 ( .x(n258), .a(B[9]), .b(A[9]) );
	aoai211_1 U81 ( .x(n236), .a(n258), .b(n278), .c(n63), .d(n193) );
	or3i_1 U82 ( .x(n182), .a(n183), .b(A[16]), .c(A[17]) );
	nor2i_1 U83 ( .x(n92), .a(n123), .b(n85) );
	inv_0 U84 ( .x(n123), .a(A[20]) );
	inv_2 U85 ( .x(n85), .a(n90) );
	nor2_1 U86 ( .x(n142), .a(n143), .b(n126) );
	inv_2 U87 ( .x(n143), .a(n189) );
	nand2i_0 U88 ( .x(n275), .a(B[14]), .b(A[14]) );
	nand2i_0 U89 ( .x(n224), .a(B[13]), .b(A[13]) );
	oai21_1 U9 ( .x(n227), .a(n61), .b(A[11]), .c(n190) );
	aoai211_1 U90 ( .x(n165), .a(n186), .b(n277), .c(n145), .d(n224) );
	inv_2 U91 ( .x(n145), .a(n188) );
	nor2_1 U92 ( .x(n144), .a(n145), .b(n125) );
	inv_2 U93 ( .x(n147), .a(n140) );
	inv_2 U94 ( .x(n229), .a(n225) );
	oai21_1 U95 ( .x(n137), .a(n155), .b(n196), .c(n229) );
	inv_2 U96 ( .x(n139), .a(n136) );
	oaoi211_1 U97 ( .x(n138), .a(n139), .b(n137), .c(n140), .d(n141) );
	nand2_2 U99 ( .x(n167), .a(n240), .b(n193) );

endmodule


module EX_test_1_desync (  ALU_result, reg_out_B_EX, mem_write_EX, mem_read_EX,
	mem_to_reg_EX, reg_write_EX, reset, IR_opcode_field, IR_function_field,
	reg_out_A, reg_out_B, Imm, reg_dst, reg_write, mem_to_reg, mem_read, mem_write,
	_byte, word, counter, test_si, test_so, test_se, sync_sel, global_g1,
	global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );

input  reset, reg_dst, reg_write, mem_to_reg, mem_read, mem_write, test_si,
	test_se, sync_sel, global_g1, global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
input [1:0] counter;
input [31:0] reg_out_A, reg_out_B, Imm;
input [5:0] IR_opcode_field, IR_function_field;
output  mem_write_EX, mem_read_EX, mem_to_reg_EX, reg_write_EX, _byte, word,
	test_so;
output [31:0] ALU_result, reg_out_B_EX;

wire ALU_result_reg_0__m2s, ALU_result_reg_10__m2s, ALU_result_reg_11__m2s,
	ALU_result_reg_12__m2s, ALU_result_reg_13__m2s, ALU_result_reg_14__m2s,
	ALU_result_reg_15__m2s, ALU_result_reg_16__m2s, ALU_result_reg_17__m2s,
	ALU_result_reg_18__m2s, ALU_result_reg_19__m2s, ALU_result_reg_1__m2s,
	ALU_result_reg_20__m2s, ALU_result_reg_21__m2s, ALU_result_reg_22__m2s,
	ALU_result_reg_23__m2s, ALU_result_reg_24__m2s, ALU_result_reg_25__m2s,
	ALU_result_reg_26__m2s, ALU_result_reg_27__m2s, ALU_result_reg_28__m2s,
	ALU_result_reg_29__m2s, ALU_result_reg_2__m2s, ALU_result_reg_30__m2s,
	ALU_result_reg_31__m2s, ALU_result_reg_3__m2s, ALU_result_reg_4__m2s,
	ALU_result_reg_5__m2s, ALU_result_reg_6__m2s, ALU_result_reg_7__m2s, ALU_result_reg_8__m2s,
	ALU_result_reg_9__m2s, N1392, N1402, N1407, N144, N1632, N1633, N1634,
	N1635, N1636, N1637, N1638, N1639, N1640, N1641, N1642, N1643, N1644,
	N1645, N1646, N1647, N1648, N1649, N1650, N1651, N1652, N1653, N1654,
	N1655, N1656, N1657, N1658, N1659, N1660, N1661, N1662, N1663, N1698,
	N1699, N1700, N1701, N1702, N1703, N1704, N1705, N1706, N1707, N1708,
	N1709, N1710, N1711, N1712, N1713, N1714, N1715, N1716, N1717, N1718,
	N1719, N1720, N1721, N1722, N1723, N1724, N1725, N1726, N1727, N1728,
	N1729, N1731, N1732, N1733, N1734, N1735, N1736, N1737, N1738, N1739,
	N1740, N1741, N1742, N1743, N1744, N1745, N1746, N1747, N1748, N1749,
	N1750, N1751, N1752, N1753, N1754, N1755, N1756, N1757, N1758, N1759,
	N1760, N1761, N1762, N1797, N1798, N1799, N1800, N1801, N1802, N1803,
	N1804, N1805, N1806, N1807, N1808, N1809, N1810, N1811, N1812, N1813,
	N1814, N1815, N1816, N1817, N1818, N1819, N1820, N1821, N1822, N1823,
	N1824, N1825, N1826, N1827, N1828, N1830, N1831, N1832, N1833, N1834,
	N1835, N1836, N1837, N1838, N1839, N1840, N1841, N1842, N1843, N1844,
	N1845, N1846, N1847, N1848, N1849, N1850, N1851, N1852, N1853, N1854,
	N1855, N1856, N1857, N1858, N1859, N1860, N1861, N1863, N1864, N1865,
	N1866, N1867, N1868, N1869, N1870, N1871, N1872, N1873, N1874, N1875,
	N1876, N1877, N1878, N1879, N1880, N1881, N1882, N1883, N1884, N1885,
	N1886, N1887, N1888, N1889, N1890, N1891, N1892, N1893, N1894, N1930,
	N1931, N1932, N1933, N1934, N1935, N1936, N1937, N1938, N1939, N1940,
	N1941, N1942, N1943, N1944, N1945, N1946, N1947, N1948, N1949, N1950,
	N1951, N1952, N1953, N1954, N1955, N1956, N1957, N1958, N1959, N1960,
	N1961, N1963, N1964, N1965, N1966, N1967, N1968, N1969, N1970, N1971,
	N1972, N1973, N1974, N1975, N1976, N1977, N1978, N1979, N1980, N1981,
	N1982, N1983, N1984, N1985, N1986, N1987, N1988, N1989, N1990, N1991,
	N1992, N1993, N1994, N1996, N1997, N1998, N1999, N2000, N2001, N2002,
	N2003, N2004, N2005, N2006, N2007, N2008, N2009, N2010, N2011, N2012,
	N2013, N2014, N2015, N2016, N2017, N2018, N2019, N2020, N2021, N2022,
	N2023, N2024, N2025, N2026, N2027, N3014, N3024, N3029, N307, N308, N309,
	N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
	N322, N323, N324, N325, N326, N327, N328, N329, N3297, N330, N3304, N331,
	N332, N333, N334, N335, N336, N337, N338, N340, N341, N342, N343, N344,
	N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355, N356,
	N357, N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
	N369, N370, N371, N69, N70, _ALU_result_reg_31_net106451, ___cell__39620_net143287,
	___cell__39620_net143326, ___cell__39620_net143595, ___cell__39620_net143596,
	___cell__39620_net143597, ___cell__39620_net143598, ___cell__39620_net143653,
	___cell__39620_net143655, ___cell__39620_net143658, ___cell__39620_net143660,
	___cell__39620_net143693, ___cell__39620_net143694, ___cell__39620_net143710,
	___cell__39620_net143720, ___cell__39620_net143722, ___cell__39620_net143735,
	___cell__39620_net143767, ___cell__39620_net143784, ___cell__39620_net143785,
	___cell__39620_net143836, ___cell__39620_net143845, ___cell__39620_net143864,
	___cell__39620_net143872, ___cell__39620_net143954, ___cell__39620_net143962,
	___cell__39620_net143982, ___cell__39620_net143983, ___cell__39620_net143997,
	___cell__39620_net144029, ___cell__39620_net144062, ___cell__39620_net144166,
	___cell__39620_net144170, ___cell__39620_net144173, ___cell__39620_net144175,
	___cell__39620_net144199, ___cell__39620_net144200, ___cell__39620_net144201,
	___cell__39620_net144257, ___cell__39620_net144302, ___cell__39620_net144303,
	___cell__39620_net144307, ___cell__39620_net144309, ___cell__39620_net144312,
	___cell__39620_net144317, ___cell__39620_net144321, ___cell__39620_net144322,
	___cell__39620_net144324, ___cell__39620_net144326, ___cell__39620_net144328,
	___cell__39620_net144329, ___cell__39620_net144330, ___cell__39620_net144331,
	___cell__39620_net144340, ___cell__39620_net144343, ___cell__39620_net144344,
	___cell__39620_net144345, ___cell__39620_net144347, ___cell__39620_net144350,
	___cell__39620_net144355, ___cell__39620_net144356, ___cell__39620_net144360,
	___cell__39620_net144374, ___cell__39620_net144406, ___cell__39620_net144517,
	___cell__39620_net144555, ___cell__39620_net144572, ___cell__39620_net144605,
	___cell__39620_net144655, ___cell__39620_net144707, ___cell__39620_net144765,
	___cell__39620_net144781, ___cell__39620_net145037, ___cell__39620_net145077,
	___cell__39620_net145078, ___cell__39620_net145150, ___cell__39620_net145190,
	___cell__39620_net145285, ___cell__39620_net145418, ___cell__39620_net145419,
	___cell__39620_net145421, ___cell__39620_net145425, ___cell__39620_net145426,
	___cell__39620_net145427, ___cell__39620_net145428, ___cell__39620_net145429,
	___cell__39620_net145444, ___cell__39620_net145450, ___cell__39620_net145451,
	___cell__39620_net145470, ___cell__39620_net145472, ___cell__39620_net145508,
	___cell__39620_net145524, ___cell__39620_net145617, ___cell__39620_net146131,
	___cell__39620_net146132, ___cell__39620_net147270, ___cell__39620_net147278,
	___cell__39620_net147296, ___cell__39620_net147350, ___cell__39620_net147731,
	___cell__39620_net147732, ___cell__39620_net147791, ___cell__6067_net21981,
	byte_reg__m2s, mem_read_EX_reg__m2s, mem_to_reg_EX_reg__m2s, mem_write_EX_reg__m2s,
	n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
	n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
	n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
	n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
	n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
	n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
	n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
	n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
	n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
	n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
	n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
	n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
	n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
	n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
	n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
	n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
	n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
	n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
	n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
	n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
	n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
	n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
	n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
	n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
	n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
	n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
	n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
	n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
	n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
	n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
	n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
	n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
	n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
	n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
	n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
	n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
	n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
	n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
	n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
	n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
	n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
	n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
	n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
	n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
	n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
	n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
	n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
	n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
	n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
	n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
	n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
	n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
	n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
	n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
	n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
	n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
	n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
	n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
	n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
	n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
	n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
	n1610, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
	n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
	n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
	n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
	n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
	n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
	n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
	n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
	n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
	n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
	n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
	n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
	n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
	n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
	n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
	n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
	n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
	n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
	n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
	n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
	n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
	n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
	n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
	n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
	n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
	n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
	n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
	n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
	n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
	n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
	n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
	n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
	n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
	n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
	n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
	n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
	n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
	n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
	n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
	n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
	n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
	n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
	n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
	n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
	n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
	n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
	n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
	n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
	n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
	n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
	n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
	n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
	n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
	n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
	n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
	n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
	n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
	n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
	n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
	n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
	n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
	n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
	n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
	n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
	n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
	n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
	n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
	n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
	n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
	n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
	n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
	n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
	n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
	n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
	n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
	n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
	n2371, n2372, n2373, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
	n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
	n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
	n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
	n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
	n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
	n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
	n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
	n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
	n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
	n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
	n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
	n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
	n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
	n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
	n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
	n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
	n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
	n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
	n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
	n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
	n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
	n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
	n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
	n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
	n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
	n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
	n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
	n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
	n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
	n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
	n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
	n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
	n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
	n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
	n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
	n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
	n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
	n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
	n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
	n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
	n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
	n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
	n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
	n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
	n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
	n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
	n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
	n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
	n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
	n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
	n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
	n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2901, n2902,
	n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
	n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
	n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
	n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
	n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
	n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
	n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
	n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
	n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
	n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
	n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
	n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
	n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
	n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
	n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
	n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
	n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
	n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
	n3083, n3084, n3085, n3086, n3088, n3089, n3090, n3091, n3092, n3093,
	n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
	n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
	n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
	n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
	n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
	n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
	n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
	n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
	n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
	n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
	n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
	n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
	n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
	n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
	n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
	n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
	n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
	n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
	n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
	n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
	n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
	n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
	n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
	n3324, n3325, n3326, n3327, n3328, n3329, n3331, n3332, n3333, n3334,
	n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
	n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
	n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
	n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
	n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
	n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
	n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
	n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
	n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
	n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
	n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
	n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
	n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465,
	n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475,
	n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
	n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
	n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505,
	n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515,
	n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525,
	n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535,
	n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545,
	n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555,
	n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565,
	n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575,
	n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585,
	n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595,
	n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605,
	n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615,
	n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625,
	n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635,
	n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645,
	n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655,
	n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665,
	n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675,
	n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685,
	n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
	n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
	n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
	n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725,
	n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735,
	n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745,
	n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755,
	n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765,
	n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775,
	n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785,
	n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795,
	n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805,
	n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815,
	n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825,
	n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835,
	n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845,
	n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855,
	n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
	n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875,
	n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885,
	n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895,
	n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905,
	n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915,
	n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925,
	n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935,
	n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945,
	n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955,
	n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965,
	n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975,
	n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
	n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
	n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
	n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015,
	n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
	n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
	n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
	n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
	n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
	n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
	n4076, n4077, n4078, n4079, n4080, n4116, n4117, n4118, n4119, n4120,
	n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
	n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
	n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4150, n4151, n4152,
	n4153, n4154, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
	n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
	n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
	n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
	n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
	n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
	n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
	n4224, n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
	n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
	n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
	n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
	n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553,
	n554, n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
	n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576, n577,
	n578, n579, n580, n581, n582, n583, n584, n585, n586, n587, n588, n589,
	n590, n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
	n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
	n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624, n625,
	n626, n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
	n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
	n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
	n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
	n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684, n685,
	n686, n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
	n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708, n709,
	n710, n711, n712, n713, n714, n715, n716, n717, n718, n719, n720, n721,
	n722, n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
	n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
	n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756, n757,
	n758, n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
	n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n782,
	n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
	n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806,
	n807, n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
	n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
	n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842,
	n843, n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
	n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
	n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878,
	n879, n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
	n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
	n903, n904, n905, n907, n908, n909, n910, n911, n912, n913, n914, n915,
	n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927,
	n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
	n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
	n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
	n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
	n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
	n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
	net149106, net149107, net149120, net149121, net149122, net149167, net149616,
	net149617, net149627, net149628, net150405, net150620, net150643, net150830,
	net151497, net151577, net151578, net151622, net151904, net152465, net156024,
	net156025, net156363, reg_out_B_EX_reg_0__m2s, reg_out_B_EX_reg_10__m2s,
	reg_out_B_EX_reg_11__m2s, reg_out_B_EX_reg_12__m2s, reg_out_B_EX_reg_13__m2s,
	reg_out_B_EX_reg_14__m2s, reg_out_B_EX_reg_15__m2s, reg_out_B_EX_reg_16__m2s,
	reg_out_B_EX_reg_17__m2s, reg_out_B_EX_reg_18__m2s, reg_out_B_EX_reg_19__m2s,
	reg_out_B_EX_reg_1__m2s, reg_out_B_EX_reg_20__m2s, reg_out_B_EX_reg_21__m2s,
	reg_out_B_EX_reg_22__m2s, reg_out_B_EX_reg_23__m2s, reg_out_B_EX_reg_24__m2s,
	reg_out_B_EX_reg_25__m2s, reg_out_B_EX_reg_26__m2s, reg_out_B_EX_reg_27__m2s,
	reg_out_B_EX_reg_28__m2s, reg_out_B_EX_reg_29__m2s, reg_out_B_EX_reg_2__m2s,
	reg_out_B_EX_reg_30__m2s, reg_out_B_EX_reg_31__m2s, reg_out_B_EX_reg_3__m2s,
	reg_out_B_EX_reg_4__m2s, reg_out_B_EX_reg_5__m2s, reg_out_B_EX_reg_6__m2s,
	reg_out_B_EX_reg_7__m2s, reg_out_B_EX_reg_8__m2s, reg_out_B_EX_reg_9__m2s,
	reg_write_EX_reg__m2s, word_reg__m2s;

	assign test_so = word;

	smlatnr_2 ALU_result_reg_0__master ( .q(ALU_result_reg_0__m2s), .qb(),
		.d(n4049), .sdi(test_si), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 ALU_result_reg_0__slave ( .q(ALU_result[0]), .qb(n4018), .d(ALU_result_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_10__master ( .q(ALU_result_reg_10__m2s), .qb(),
		.d(n4059), .sdi(ALU_result[9]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_10__slave ( .q(ALU_result[10]), .qb(n4020), .d(ALU_result_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 ALU_result_reg_11__master ( .q(ALU_result_reg_11__m2s), .qb(),
		.d(n4060), .sdi(ALU_result[10]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 ALU_result_reg_11__slave ( .q(ALU_result[11]), .qb(n4021), .d(ALU_result_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_12__master ( .q(ALU_result_reg_12__m2s), .qb(),
		.d(n4061), .sdi(ALU_result[11]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_12__slave ( .q(ALU_result[12]), .qb(n4154), .d(ALU_result_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_13__master ( .q(ALU_result_reg_13__m2s), .qb(),
		.d(n4062), .sdi(n4154), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_13__slave ( .q(ALU_result[13]), .qb(n4022), .d(ALU_result_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_14__master ( .q(ALU_result_reg_14__m2s), .qb(),
		.d(n4063), .sdi(ALU_result[13]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_14__slave ( .q(ALU_result[14]), .qb(n4153), .d(ALU_result_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_15__master ( .q(ALU_result_reg_15__m2s), .qb(),
		.d(n4064), .sdi(n4153), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_15__slave ( .q(ALU_result[15]), .qb(n4023), .d(ALU_result_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_16__master ( .q(ALU_result_reg_16__m2s), .qb(),
		.d(n4065), .sdi(ALU_result[15]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_16__slave ( .q(ALU_result[16]), .qb(n4024), .d(ALU_result_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_17__master ( .q(ALU_result_reg_17__m2s), .qb(),
		.d(n4066), .sdi(ALU_result[16]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_17__slave ( .q(ALU_result[17]), .qb(n4025), .d(ALU_result_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_18__master ( .q(ALU_result_reg_18__m2s), .qb(),
		.d(n4067), .sdi(ALU_result[17]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_18__slave ( .q(ALU_result[18]), .qb(n4152), .d(ALU_result_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_19__master ( .q(ALU_result_reg_19__m2s), .qb(),
		.d(n4068), .sdi(n4152), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_19__slave ( .q(ALU_result[19]), .qb(n4151), .d(ALU_result_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_1__master ( .q(ALU_result_reg_1__m2s), .qb(),
		.d(n4050), .sdi(ALU_result[0]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_1__slave ( .q(ALU_result[1]), .qb(n4019), .d(ALU_result_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 ALU_result_reg_20__master ( .q(ALU_result_reg_20__m2s), .qb(),
		.d(n4069), .sdi(n4151), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 ALU_result_reg_20__slave ( .q(ALU_result[20]), .qb(n4027), .d(ALU_result_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_21__master ( .q(ALU_result_reg_21__m2s), .qb(),
		.d(n4070), .sdi(ALU_result[20]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_21__slave ( .q(ALU_result[21]), .qb(n4028), .d(ALU_result_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_22__master ( .q(ALU_result_reg_22__m2s), .qb(),
		.d(n4071), .sdi(ALU_result[21]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_22__slave ( .q(ALU_result[22]), .qb(n4029), .d(ALU_result_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_23__master ( .q(ALU_result_reg_23__m2s), .qb(),
		.d(n4072), .sdi(ALU_result[22]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_23__slave ( .q(ALU_result[23]), .qb(n4030), .d(ALU_result_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_24__master ( .q(ALU_result_reg_24__m2s), .qb(),
		.d(n4073), .sdi(ALU_result[23]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_24__slave ( .q(ALU_result[24]), .qb(n4031), .d(ALU_result_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_25__master ( .q(ALU_result_reg_25__m2s), .qb(),
		.d(n4074), .sdi(ALU_result[24]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_25__slave ( .q(ALU_result[25]), .qb(n4032), .d(ALU_result_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_26__master ( .q(ALU_result_reg_26__m2s), .qb(),
		.d(n4075), .sdi(ALU_result[25]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_26__slave ( .q(ALU_result[26]), .qb(n4033), .d(ALU_result_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_27__master ( .q(ALU_result_reg_27__m2s), .qb(),
		.d(n4076), .sdi(ALU_result[26]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_27__slave ( .q(ALU_result[27]), .qb(n4034), .d(ALU_result_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_28__master ( .q(ALU_result_reg_28__m2s), .qb(),
		.d(n4077), .sdi(ALU_result[27]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_28__slave ( .q(ALU_result[28]), .qb(n4035), .d(ALU_result_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 ALU_result_reg_29__master ( .q(ALU_result_reg_29__m2s), .qb(),
		.d(n4078), .sdi(ALU_result[28]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 ALU_result_reg_29__slave ( .q(ALU_result[29]), .qb(n4036), .d(ALU_result_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_2__master ( .q(ALU_result_reg_2__m2s), .qb(),
		.d(n4051), .sdi(ALU_result[1]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_2__slave ( .q(ALU_result[2]), .qb(n4026), .d(ALU_result_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 ALU_result_reg_30__master ( .q(ALU_result_reg_30__m2s), .qb(),
		.d(n4079), .sdi(ALU_result[29]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 ALU_result_reg_30__slave ( .q(ALU_result[30]), .qb(n4038), .d(ALU_result_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 ALU_result_reg_31__master ( .q(ALU_result_reg_31__m2s), .qb(),
		.d(_ALU_result_reg_31_net106451), .sdi(ALU_result[30]), .se(test_se),
		.g(Ctrl__Regs_1__en1), .rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 ALU_result_reg_31__slave ( .q(ALU_result[31]), .qb(n4039), .d(ALU_result_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_3__master ( .q(ALU_result_reg_3__m2s), .qb(),
		.d(n4052), .sdi(ALU_result[2]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_3__slave ( .q(ALU_result[3]), .qb(n4037), .d(ALU_result_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_4__master ( .q(ALU_result_reg_4__m2s), .qb(),
		.d(n4053), .sdi(ALU_result[3]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_4__slave ( .q(ALU_result[4]), .qb(n4040), .d(ALU_result_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_5__master ( .q(ALU_result_reg_5__m2s), .qb(),
		.d(n4054), .sdi(ALU_result[4]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4017), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_5__slave ( .q(ALU_result[5]), .qb(n4041), .d(ALU_result_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_6__master ( .q(ALU_result_reg_6__m2s), .qb(),
		.d(n4055), .sdi(ALU_result[5]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_6__slave ( .q(ALU_result[6]), .qb(n4042), .d(ALU_result_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_7__master ( .q(ALU_result_reg_7__m2s), .qb(),
		.d(n4056), .sdi(ALU_result[6]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 ALU_result_reg_7__slave ( .q(ALU_result[7]), .qb(n4043), .d(ALU_result_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_8__master ( .q(ALU_result_reg_8__m2s), .qb(),
		.d(n4057), .sdi(ALU_result[7]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 ALU_result_reg_8__slave ( .q(ALU_result[8]), .qb(n4044), .d(ALU_result_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 ALU_result_reg_9__master ( .q(ALU_result_reg_9__m2s), .qb(),
		.d(n4058), .sdi(ALU_result[8]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n543), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 ALU_result_reg_9__slave ( .q(ALU_result[9]), .qb(n4045), .d(ALU_result_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	oai21_1 U100 ( .x(n3235), .a(n1577), .b(n1729), .c(n665) );
	inv_2 U1000 ( .x(n1964), .a(n1070) );
	nor2i_0 U1001 ( .x(n1235), .a(Imm[7]), .b(n734) );
	aoi21_1 U1002 ( .x(n2635), .a(N1754), .b(___cell__39620_net145150), .c(n1235) );
	nand2i_2 U1003 ( .x(n2639), .a(n1801), .b(n809) );
	inv_2 U1004 ( .x(n1801), .a(N1655) );
	nand2_2 U1005 ( .x(n2631), .a(n829), .b(n634) );
	nand2i_2 U1006 ( .x(n2638), .a(n2631), .b(___cell__39620_net145285) );
	nand2i_2 U1007 ( .x(n2645), .a(n1805), .b(n1987) );
	inv_2 U1008 ( .x(n1805), .a(N1820) );
	inv_5 U1009 ( .x(n1315), .a(n2722) );
	ao21_1 U101 ( .x(n3236), .a(n1147), .b(n1136), .c(n3235) );
	nand2i_2 U1010 ( .x(n2644), .a(n1055), .b(n2557) );
	inv_2 U1011 ( .x(n661), .a(n869) );
	inv_5 U1012 ( .x(n3648), .a(n844) );
	inv_2 U1013 ( .x(n1804), .a(N1953) );
	nand2i_2 U1014 ( .x(___cell__39620_net143845), .a(___cell__39620_net144360),
		.b(n708) );
	nor2i_1 U1015 ( .x(n1236), .a(N1986), .b(___cell__39620_net143845) );
	oai211_2 U1016 ( .x(n3821), .a(n3460), .b(n1623), .c(n2602), .d(n3820) );
	nor2i_3 U1017 ( .x(n1233), .a(___cell__39620_net143864), .b(n1234) );
	inv_8 U1018 ( .x(n1322), .a(n1972) );
	oai221_4 U1019 ( .x(n2609), .a(n3418), .b(n4004), .c(n1322), .d(n1565),
		.e(n1807) );
	nand2i_2 U102 ( .x(n3234), .a(n1625), .b(n2806) );
	aoi22_1 U1020 ( .x(n2608), .a(n649), .b(n2609), .c(n650), .d(n2574) );
	oai21_1 U1021 ( .x(n2604), .a(n1486), .b(n690), .c(n2605) );
	inv_2 U1022 ( .x(n1063), .a(n646) );
	inv_2 U1023 ( .x(n2607), .a(n3826) );
	nand2i_0 U1024 ( .x(n2620), .a(___cell__39620_net144707), .b(___cell__39620_net145617) );
	inv_8 U1025 ( .x(n811), .a(n606) );
	nor2i_1 U1026 ( .x(n1228), .a(N1854), .b(n946) );
	inv_2 U1027 ( .x(n1230), .a(N1821) );
	nor2_1 U1028 ( .x(n1229), .a(n1077), .b(n1230) );
	inv_2 U1029 ( .x(n1795), .a(N1954) );
	mux2i_1 U103 ( .x(n3239), .d0(___cell__39620_net144201), .sl(net152465),
		.d1(___cell__39620_net145285) );
	inv_2 U1030 ( .x(n1794), .a(N1887) );
	nand2i_2 U1031 ( .x(n2595), .a(n1794), .b(n3997) );
	nor2i_1 U1032 ( .x(n1226), .a(N1755), .b(___cell__39620_net143710) );
	aoi211_1 U1033 ( .x(n2594), .a(N1722), .b(___cell__39620_net145190), .c(n1227),
		.d(n1226) );
	nand2i_2 U1034 ( .x(n2593), .a(n1793), .b(n809) );
	inv_2 U1035 ( .x(n1793), .a(N1656) );
	inv_2 U1036 ( .x(n1788), .a(N1955) );
	inv_2 U1037 ( .x(n1214), .a(N1822) );
	nor2_1 U1038 ( .x(n1213), .a(n1077), .b(n1214) );
	oai221_3 U1039 ( .x(n565), .a(n1302), .b(n1043), .c(n3524), .d(n4007),
		.e(n1806) );
	nand2i_2 U104 ( .x(n1653), .a(n497), .b(n676) );
	aoi21_1 U1040 ( .x(n2546), .a(N1756), .b(___cell__39620_net145150), .c(n1212) );
	nand2i_2 U1041 ( .x(n2549), .a(n1785), .b(n809) );
	inv_2 U1042 ( .x(n1785), .a(N1657) );
	nand2_2 U1043 ( .x(n2545), .a(n689), .b(n590) );
	nand2i_2 U1044 ( .x(n2548), .a(n2545), .b(___cell__39620_net145285) );
	nor2_1 U1045 ( .x(n1060), .a(n1061), .b(n645) );
	nand2i_2 U1046 ( .x(n1531), .a(IR_function_field[1]), .b(IR_function_field[0]) );
	aoi21_1 U1047 ( .x(n2566), .a(___cell__39620_net144517), .b(n2375), .c(n2564) );
	nand2i_2 U1048 ( .x(n3811), .a(n1625), .b(n2649) );
	inv_5 U1049 ( .x(n2266), .a(n1091) );
	nor2_1 U105 ( .x(n1427), .a(n1428), .b(n1429) );
	nand3_1 U1050 ( .x(n3812), .a(n2562), .b(n3811), .c(n2566) );
	nand2i_2 U1051 ( .x(n2584), .a(n688), .b(___cell__39620_net145617) );
	inv_8 U1052 ( .x(n3385), .a(n3384) );
	inv_2 U1053 ( .x(n3444), .a(n3443) );
	nor2i_1 U1054 ( .x(n1650), .a(n2001), .b(n1539) );
	oai22_1 U1055 ( .x(n2560), .a(n2475), .b(n1687), .c(n1648), .d(n1690) );
	aoi21_1 U1056 ( .x(n2561), .a(n1256), .b(n2477), .c(n2560) );
	nand2i_2 U1057 ( .x(n3815), .a(n1578), .b(n3684) );
	inv_5 U1058 ( .x(n1578), .a(reg_out_A[24]) );
	inv_2 U1059 ( .x(n3447), .a(n2738) );
	nor2_1 U106 ( .x(n3232), .a(n3229), .b(n3230) );
	nand2_2 U1060 ( .x(n3813), .a(n1249), .b(n2738) );
	nor2i_1 U1061 ( .x(n1220), .a(n1221), .b(n1222) );
	inv_2 U1062 ( .x(n1222), .a(n2492) );
	nand2i_2 U1063 ( .x(n2572), .a(n1484), .b(n2139) );
	exnor2_1 U1064 ( .x(n1483), .a(n590), .b(n689) );
	oai21_1 U1065 ( .x(n2571), .a(n1483), .b(n690), .c(n2572) );
	nor2_0 U1066 ( .x(n2543), .a(n1626), .b(net149120) );
	nand2i_2 U1067 ( .x(n1218), .a(n1781), .b(n530) );
	aoi21_1 U1068 ( .x(n1216), .a(n1217), .b(n1218), .c(n1219) );
	nor2i_1 U1069 ( .x(n2544), .a(n1451), .b(n670) );
	nor2_1 U107 ( .x(n3228), .a(n3226), .b(n3227) );
	nand4_1 U1070 ( .x(n3782), .a(n2480), .b(n3781), .c(n2479), .d(n3780) );
	inv_2 U1071 ( .x(n2435), .a(n1711) );
	inv_2 U1072 ( .x(n2436), .a(n1712) );
	nand2i_2 U1073 ( .x(n3780), .a(n1623), .b(n2649) );
	nand2i_2 U1074 ( .x(n1443), .a(n1659), .b(n1542) );
	inv_2 U1075 ( .x(n1542), .a(n1539) );
	nand2i_2 U1076 ( .x(n1539), .a(IR_function_field[5]), .b(n1540) );
	inv_2 U1077 ( .x(n1540), .a(n1538) );
	inv_2 U1078 ( .x(n1661), .a(n1443) );
	oai22_1 U1079 ( .x(n2474), .a(n1648), .b(n1715), .c(n2475), .d(n1713) );
	nor2_1 U108 ( .x(n3225), .a(n3223), .b(n3224) );
	aoi21_1 U1080 ( .x(n2476), .a(n1249), .b(n2477), .c(n2474) );
	nand2i_2 U1081 ( .x(n3784), .a(n4009), .b(n2286) );
	oai211_2 U1082 ( .x(n2286), .a(n507), .b(n1546), .c(n3407), .d(n3408) );
	aoi21_1 U1083 ( .x(n2478), .a(n1256), .b(n2373), .c(n1194) );
	nand2i_2 U1084 ( .x(___cell__39620_net144302), .a(n1533), .b(n675) );
	nor2i_0 U1085 ( .x(n1619), .a(IR_opcode_field[0]), .b(n1519) );
	nand2_2 U1086 ( .x(n1618), .a(n1619), .b(___cell__39620_net144303) );
	inv_2 U1087 ( .x(n1061), .a(n1531) );
	nand2i_2 U1088 ( .x(n1525), .a(n1523), .b(n1526) );
	nand2_2 U1089 ( .x(n3798), .a(n1249), .b(n2779) );
	nor2_1 U109 ( .x(n3222), .a(n3220), .b(n3221) );
	inv_2 U1090 ( .x(n3684), .a(n1093) );
	nand2i_2 U1091 ( .x(n3799), .a(n1219), .b(n3684) );
	nand2_2 U1092 ( .x(n3797), .a(n1714), .b(n2306) );
	inv_2 U1093 ( .x(n1150), .a(n1687) );
	aoi222_1 U1094 ( .x(n2518), .a(n1256), .b(n2433), .c(n1150), .d(n2270),
		.e(n2273), .f(n904) );
	nand2i_2 U1095 ( .x(n1590), .a(IR_function_field[2]), .b(n1526) );
	inv_2 U1096 ( .x(n1526), .a(n1522) );
	or3i_1 U1097 ( .x(n1522), .a(IR_function_field[5]), .b(IR_function_field[4]),
		.c(IR_function_field[3]) );
	inv_8 U1098 ( .x(n1217), .a(n1700) );
	inv_5 U1099 ( .x(n3779), .a(n3778) );
	nor2_1 U110 ( .x(n3281), .a(n1939), .b(n1951) );
	nand2i_2 U1100 ( .x(n3806), .a(n670), .b(n3778) );
	inv_14 U1101 ( .x(n915), .a(n813) );
	inv_2 U1102 ( .x(n3386), .a(n2568) );
	exnor2_1 U1103 ( .x(n1481), .a(n540), .b(Imm[26]) );
	inv_2 U1104 ( .x(n3810), .a(n1481) );
	inv_2 U1105 ( .x(___cell__39620_net144201), .a(___cell__39620_net144199) );
	nand2_2 U1106 ( .x(n1116), .a(___cell__39620_net147732), .b(___cell__39620_net144201) );
	nand2_2 U1107 ( .x(n2526), .a(n2193), .b(n3810) );
	exnor2_1 U1108 ( .x(n1482), .a(n540), .b(reg_out_B[26]) );
	nand2i_2 U1109 ( .x(n2525), .a(n1482), .b(n2139) );
	inv_5 U111 ( .x(n1093), .a(n737) );
	nand2_2 U1110 ( .x(n3801), .a(n3315), .b(n855) );
	inv_10 U1111 ( .x(n882), .a(n825) );
	inv_2 U1112 ( .x(n2432), .a(n1122) );
	oai21_1 U1113 ( .x(n3739), .a(n536), .b(n3738), .c(n1807) );
	inv_2 U1114 ( .x(n3738), .a(n2629) );
	inv_2 U1115 ( .x(n854), .a(n1807) );
	inv_2 U1116 ( .x(n1330), .a(n1565) );
	nand2i_4 U1117 ( .x(n2981), .a(n3585), .b(n3783) );
	nand2i_2 U1118 ( .x(n3425), .a(n1565), .b(n2981) );
	nand2i_0 U1119 ( .x(n3424), .a(n1559), .b(n1728) );
	nor2i_1 U112 ( .x(n1442), .a(n1443), .b(n1444) );
	nand2i_2 U1120 ( .x(n1582), .a(n1451), .b(n1545) );
	nand2_2 U1121 ( .x(n3762), .a(n3343), .b(n855) );
	nand2i_2 U1124 ( .x(n1160), .a(n1568), .b(n1543) );
	nor2i_1 U1125 ( .x(n1612), .a(IR_opcode_field[0]), .b(IR_opcode_field[1]) );
	inv_8 U1126 ( .x(n1302), .a(n2677) );
	nor2_1 U1127 ( .x(n1207), .a(n734), .b(n1208) );
	nand2i_3 U1128 ( .x(n2506), .a(n1775), .b(n809) );
	nand2_0 U1129 ( .x(n2502), .a(Imm[26]), .b(n540) );
	oai21_1 U113 ( .x(n3280), .a(n1442), .b(n1093), .c(n3281) );
	nand2i_2 U1130 ( .x(n2505), .a(n2502), .b(___cell__39620_net147791) );
	nand2i_2 U1131 ( .x(___cell__39620_net144360), .a(n675), .b(n810) );
	oai21_3 U1132 ( .x(n3726), .a(n4125), .b(n1290), .c(n1806) );
	inv_8 U1133 ( .x(n1198), .a(n2423) );
	nand2i_2 U1134 ( .x(n2363), .a(n1742), .b(n2837) );
	inv_2 U1135 ( .x(n1742), .a(N310) );
	inv_2 U1136 ( .x(n571), .a(n3435) );
	nand2i_1 U1137 ( .x(n2361), .a(n1186), .b(n2197) );
	nand2i_2 U1138 ( .x(n2356), .a(n621), .b(n3757) );
	oai21_1 U1139 ( .x(n2352), .a(n1473), .b(n690), .c(n2353) );
	nor2_1 U114 ( .x(n3275), .a(n3272), .b(n3273) );
	nand4i_1 U1140 ( .x(n2354), .a(n2352), .b(n2355), .c(n2356), .d(n2357) );
	inv_2 U1141 ( .x(___cell__39620_net145524), .a(___cell__39620_net145444) );
	oai221_1 U1142 ( .x(n2365), .a(n2366), .b(n1647), .c(___cell__39620_net145524),
		.d(n1646), .e(n2367) );
	nand4i_1 U1143 ( .x(n2364), .a(n2365), .b(n2368), .c(n2369), .d(n2370) );
	nand4_1 U1144 ( .x(n1173), .a(n2347), .b(n2345), .c(n2348), .d(n2349) );
	nand2i_2 U1145 ( .x(n2347), .a(n1182), .b(n2168) );
	nand2i_2 U1146 ( .x(n2348), .a(n1055), .b(n2165) );
	nand2i_2 U1147 ( .x(n2349), .a(n1743), .b(n809) );
	inv_2 U1148 ( .x(n1743), .a(N1635) );
	nor2i_1 U1149 ( .x(n1167), .a(N1833), .b(n946) );
	and3i_1 U115 ( .x(n3271), .a(n3264), .b(n3265), .c(n3268) );
	nor2i_1 U1150 ( .x(n1168), .a(N1999), .b(n1169) );
	aoi211_1 U1151 ( .x(n1172), .a(N1966), .b(___cell__39620_net145508), .c(n1168),
		.d(n1167) );
	inv_2 U1152 ( .x(n1745), .a(N1933) );
	nand2i_2 U1153 ( .x(n1171), .a(n1745), .b(n3662) );
	nor2i_2 U1154 ( .x(n1164), .a(n1165), .b(n1166) );
	aoi21_1 U1155 ( .x(n2346), .a(N1701), .b(___cell__39620_net145190), .c(n1163) );
	inv_2 U1156 ( .x(n1746), .a(N1800) );
	nand2i_2 U1157 ( .x(n2351), .a(n1746), .b(n1987) );
	inv_2 U1158 ( .x(n1744), .a(N1866) );
	nand2i_2 U1159 ( .x(n2350), .a(n1744), .b(n3997) );
	nor2_1 U116 ( .x(n3263), .a(n3261), .b(n3262) );
	aoi221_1 U1160 ( .x(n2836), .a(n692), .b(n1733), .c(n917), .d(___cell__39620_net145444),
		.e(n2838) );
	nand2i_2 U1161 ( .x(n2835), .a(n1647), .b(n3705) );
	inv_2 U1162 ( .x(n1589), .a(n1582) );
	oai211_2 U1163 ( .x(n2834), .a(n2360), .b(n1588), .c(n2835), .d(n2836) );
	inv_5 U1164 ( .x(n1428), .a(n1639) );
	ao22_2 U1165 ( .x(n2825), .a(n502), .b(n2826), .c(n1267), .d(n2827) );
	inv_2 U1166 ( .x(n2829), .a(n1496) );
	aoi21_1 U1167 ( .x(n2828), .a(n2139), .b(n2829), .c(n1284) );
	aoai211_1 U1168 ( .x(n2824), .a(n692), .b(n530), .c(n1064), .d(n815) );
	nand2i_2 U1169 ( .x(n2823), .a(n670), .b(n3757) );
	nor3i_1 U117 ( .x(n3260), .a(n1518), .b(n3258), .c(n3259) );
	inv_2 U1170 ( .x(n1436), .a(n1620) );
	inv_2 U1171 ( .x(n2822), .a(n3760) );
	aoi211_1 U1172 ( .x(n2814), .a(N1733), .b(___cell__39620_net145150), .c(n1271),
		.d(n1270) );
	inv_2 U1173 ( .x(n1838), .a(N1634) );
	nand2i_2 U1174 ( .x(n2816), .a(n1838), .b(n809) );
	nand2i_2 U1175 ( .x(n2815), .a(n1182), .b(n2165) );
	inv_2 U1176 ( .x(n1839), .a(N1932) );
	nand2i_2 U1177 ( .x(n2820), .a(n1839), .b(n3999) );
	inv_2 U1178 ( .x(n1841), .a(N1965) );
	nand2i_2 U1179 ( .x(n2819), .a(n1841), .b(___cell__39620_net145508) );
	inv_5 U118 ( .x(n1585), .a(n608) );
	inv_2 U1180 ( .x(n1840), .a(N1832) );
	nand2i_2 U1181 ( .x(n2818), .a(n1840), .b(n4000) );
	nand2i_2 U1182 ( .x(n1275), .a(n1842), .b(n3624) );
	inv_2 U1183 ( .x(n1842), .a(N1998) );
	inv_2 U1184 ( .x(n1692), .a(N313) );
	inv_2 U1185 ( .x(n2142), .a(n2197) );
	oai211_1 U1186 ( .x(n2141), .a(n2142), .b(n1566), .c(n2138), .d(n2134) );
	nand2i_2 U1187 ( .x(n2155), .a(n621), .b(n3693) );
	aoi22_1 U1188 ( .x(n2156), .a(n2157), .b(n1085), .c(n2106), .d(n1204) );
	inv_2 U1189 ( .x(n1693), .a(N346) );
	exnor2_1 U119 ( .x(n1508), .a(reg_out_B[14]), .b(n644) );
	inv_2 U1190 ( .x(n1694), .a(N2002) );
	inv_2 U1191 ( .x(n1696), .a(N1936) );
	nand2i_2 U1192 ( .x(n3697), .a(n1696), .b(n3999) );
	inv_2 U1193 ( .x(n1699), .a(N1969) );
	nand2i_2 U1194 ( .x(n2125), .a(n1699), .b(___cell__39620_net145508) );
	inv_2 U1195 ( .x(n1698), .a(N1803) );
	nand2i_2 U1196 ( .x(n2124), .a(n1698), .b(n1987) );
	inv_2 U1197 ( .x(n1697), .a(N1836) );
	nand2i_2 U1198 ( .x(n2123), .a(n1697), .b(n4000) );
	and4i_1 U1199 ( .x(n2122), .a(n2121), .b(n2123), .c(n2124), .d(n2125) );
	nand2_2 U120 ( .x(n3631), .a(n3559), .b(___cell__39620_net144331) );
	aoi21_1 U1200 ( .x(n2120), .a(N1704), .b(___cell__39620_net145190), .c(n1111) );
	inv_2 U1201 ( .x(n1695), .a(N1638) );
	nand2i_2 U1202 ( .x(n2119), .a(n1695), .b(n809) );
	nand2i_2 U1203 ( .x(n2118), .a(n1166), .b(n2168) );
	aoi22_1 U1204 ( .x(n3104), .a(n650), .b(n3078), .c(n1221), .d(n3000) );
	aoi221_1 U1205 ( .x(n3101), .a(n1204), .b(n3075), .c(n649), .d(n2014),
		.e(n3102) );
	aoi21_1 U1206 ( .x(n3109), .a(n2022), .b(n3110), .c(n1389) );
	aoi222_1 U1207 ( .x(n3115), .a(n3118), .b(___cell__39620_net143864), .c(n894),
		.d(n1700), .e(ALU_result[12]), .f(n3057) );
	nand2i_2 U1208 ( .x(n3107), .a(n1900), .b(n977) );
	inv_2 U1209 ( .x(n1900), .a(N352) );
	nand2i_2 U121 ( .x(n3961), .a(n1625), .b(n3291) );
	inv_2 U1210 ( .x(n1906), .a(N1975) );
	nand2i_2 U1211 ( .x(n3096), .a(n1906), .b(___cell__39620_net145508) );
	inv_2 U1212 ( .x(n1905), .a(N1842) );
	nand2i_2 U1213 ( .x(n3095), .a(n1905), .b(n735) );
	aoi22_1 U1214 ( .x(n3094), .a(n1095), .b(n1988), .c(n1197), .d(n1397) );
	aoi21_1 U1215 ( .x(n3093), .a(n662), .b(n594), .c(n1381) );
	nand4_1 U1216 ( .x(n1386), .a(n3093), .b(n3094), .c(n3095), .d(n3096) );
	nand2i_2 U1217 ( .x(n1385), .a(n1901), .b(n3624) );
	inv_2 U1218 ( .x(n1901), .a(N2008) );
	inv_2 U1219 ( .x(n1904), .a(N1942) );
	ao22_2 U122 ( .x(n712), .a(n526), .b(n1256), .c(n504), .d(n3020) );
	nand2i_2 U1220 ( .x(n1384), .a(n1904), .b(n3999) );
	nor2i_3 U1221 ( .x(n1379), .a(n1380), .b(n1055) );
	inv_2 U1222 ( .x(n1903), .a(N1875) );
	nand2i_2 U1223 ( .x(n3092), .a(n1903), .b(n3997) );
	aoi211_1 U1224 ( .x(n3090), .a(N1644), .b(n809), .c(n1378), .d(n1376) );
	inv_2 U1225 ( .x(n1902), .a(N1743) );
	nand2i_2 U1226 ( .x(n3091), .a(n1902), .b(___cell__39620_net145150) );
	and4i_1 U1227 ( .x(n1383), .a(n1379), .b(n3091), .c(n3090), .d(n3092) );
	inv_2 U1228 ( .x(n1675), .a(N347) );
	nand2i_2 U1229 ( .x(n2095), .a(n1675), .b(n977) );
	nand2_2 U123 ( .x(n3547), .a(n3548), .b(n3549) );
	aoi22_1 U1231 ( .x(n2088), .a(n649), .b(n2089), .c(n650), .d(n2090) );
	nand4_1 U1232 ( .x(n2094), .a(n2091), .b(n2088), .c(n2092), .d(n2095) );
	inv_2 U1233 ( .x(n589), .a(n2135) );
	aoi221_3 U1234 ( .x(n2096), .a(n2106), .b(___cell__39620_net143864), .c(n2107),
		.d(n1204), .e(n2103) );
	inv_2 U1235 ( .x(n1681), .a(N1970) );
	nand2i_2 U1236 ( .x(n2077), .a(n1681), .b(___cell__39620_net145508) );
	inv_2 U1237 ( .x(n1680), .a(N1804) );
	nand2i_2 U1238 ( .x(n2076), .a(n1680), .b(n1987) );
	aoi22_1 U1239 ( .x(n2074), .a(n1318), .b(n1993), .c(n662), .d(n1992) );
	inv_5 U124 ( .x(n2273), .a(n1690) );
	aoi21_1 U1240 ( .x(n2075), .a(n1197), .b(n2043), .c(n1099) );
	nand4_1 U1241 ( .x(n1103), .a(n2075), .b(n2074), .c(n2076), .d(n2077) );
	nand2i_2 U1242 ( .x(n1102), .a(n1677), .b(n3624) );
	inv_2 U1243 ( .x(n1677), .a(N2003) );
	inv_2 U1244 ( .x(n1679), .a(N1937) );
	nand2i_2 U1245 ( .x(n1101), .a(n1679), .b(n3662) );
	nand2i_2 U1246 ( .x(n2071), .a(n2068), .b(___cell__39620_net145285) );
	inv_2 U1247 ( .x(n1678), .a(N1639) );
	nand2i_2 U1248 ( .x(n2072), .a(n1678), .b(n809) );
	nand2i_2 U1249 ( .x(n2501), .a(___cell__39620_net144406), .b(n3785) );
	inv_4 U125 ( .x(n3352), .a(n658) );
	nand2i_2 U1250 ( .x(n2500), .a(n784), .b(n3782) );
	aoi21_1 U1251 ( .x(n2498), .a(n1085), .b(n2499), .c(n1206) );
	nand2i_2 U1253 ( .x(n2496), .a(n1761), .b(n2837) );
	inv_2 U1254 ( .x(n1761), .a(N334) );
	and4i_3 U1255 ( .x(n2493), .a(n2494), .b(n2491), .c(n2488), .d(n2484) );
	aoi22_1 U1256 ( .x(n2491), .a(n650), .b(n2492), .c(n1221), .d(n2400) );
	aoi22_1 U1257 ( .x(n2488), .a(n539), .b(n2489), .c(n535), .d(n2490) );
	and4i_3 U1258 ( .x(n2484), .a(n2481), .b(n2485), .c(n2486), .d(n2487) );
	inv_2 U1259 ( .x(n2494), .a(n3794) );
	and2_5 U126 ( .x(n512), .a(n3352), .b(n3353) );
	nand2i_2 U1260 ( .x(n3794), .a(n1566), .b(n3422) );
	inv_5 U1261 ( .x(n1760), .a(reg_out_B[27]) );
	inv_5 U1262 ( .x(n680), .a(Imm[27]) );
	oai21_2 U1263 ( .x(n2399), .a(n3419), .b(n1565), .c(n3571) );
	aoi222_1 U1264 ( .x(n2495), .a(n1191), .b(n2399), .c(n681), .d(___cell__39620_net145617),
		.e(reg_out_B[27]), .f(n1064) );
	inv_8 U1265 ( .x(n1573), .a(reg_out_A[26]) );
	inv_2 U1266 ( .x(n1769), .a(N1857) );
	nand2i_2 U1267 ( .x(n2472), .a(n1769), .b(n735) );
	inv_2 U1268 ( .x(n1768), .a(N1824) );
	nand2i_2 U1269 ( .x(n2471), .a(n1768), .b(n1987) );
	oai22_1 U127 ( .x(n2131), .a(n512), .b(n1687), .c(n1570), .d(n1690) );
	inv_2 U1270 ( .x(n1770), .a(N1990) );
	nand2i_2 U1271 ( .x(n2470), .a(n1770), .b(___cell__39620_net145508) );
	aoi21_1 U1272 ( .x(n2469), .a(n1095), .b(n2473), .c(n1196) );
	nand2i_2 U1273 ( .x(n1201), .a(n1763), .b(n3624) );
	inv_2 U1274 ( .x(n1763), .a(N2023) );
	inv_2 U1275 ( .x(n1162), .a(n2384) );
	inv_2 U1276 ( .x(n1764), .a(N1659) );
	inv_2 U1277 ( .x(n1765), .a(N1725) );
	aoi21_1 U1278 ( .x(n3244), .a(___cell__39620_net143785), .b(n3245), .c(n1438) );
	and4i_3 U1279 ( .x(n3248), .a(n3251), .b(n3253), .c(n3254), .d(n3255) );
	nor2i_0 U128 ( .x(n1110), .a(n922), .b(n1093) );
	ao21_3 U1280 ( .x(n1440), .a(n3992), .b(n3991), .c(n1609) );
	inv_2 U1281 ( .x(n2004), .a(n1937) );
	inv_2 U1282 ( .x(n1638), .a(n1627) );
	aoi221_1 U1283 ( .x(n3290), .a(n1638), .b(n3214), .c(N340), .d(n1597),
		.e(n1445) );
	aoi221_3 U1284 ( .x(n3287), .a(n1576), .b(n3288), .c(n1589), .d(n3289),
		.e(n1453) );
	nand2i_2 U1285 ( .x(n3131), .a(n1574), .b(n2014) );
	oai21_1 U1287 ( .x(n3129), .a(n3130), .b(n1566), .c(n3131) );
	nand2i_2 U1288 ( .x(n3134), .a(n1908), .b(n2837) );
	inv_2 U1289 ( .x(n1908), .a(N318) );
	nand2i_2 U1290 ( .x(n3133), .a(n1588), .b(n3078) );
	oai211_1 U1291 ( .x(n3126), .a(n1403), .b(n1907), .c(n3127), .d(n3128) );
	aoi21_1 U1292 ( .x(n3132), .a(n1221), .b(n3041), .c(n3126) );
	nand2_1 U1293 ( .x(n3147), .a(n1085), .b(n3117) );
	nand2_2 U1294 ( .x(n3146), .a(n3170), .b(___cell__39620_net143864) );
	inv_5 U1295 ( .x(n900), .a(reg_out_A[11]) );
	nand2i_2 U1296 ( .x(n3137), .a(n1909), .b(n977) );
	inv_2 U1297 ( .x(n1909), .a(N351) );
	inv_14 U1298 ( .x(___cell__39620_net144655), .a(Imm[11]) );
	and4i_3 U1299 ( .x(n3135), .a(n3139), .b(n3141), .c(n3142), .d(n3143) );
	nand2i_2 U130 ( .x(n3710), .a(n4008), .b(n2806) );
	nand2_2 U1300 ( .x(n3141), .a(n2024), .b(n3116) );
	nand2_2 U1301 ( .x(n3142), .a(n2022), .b(n3113) );
	inv_2 U1302 ( .x(n1915), .a(N1974) );
	nand2i_2 U1303 ( .x(n3125), .a(n1915), .b(___cell__39620_net145508) );
	inv_2 U1304 ( .x(n1914), .a(N1808) );
	nand2i_2 U1305 ( .x(n3124), .a(n1914), .b(n1987) );
	aoi22_1 U1306 ( .x(n3123), .a(n1095), .b(n1054), .c(n1197), .d(n1988) );
	nand2i_2 U1307 ( .x(n1401), .a(n1910), .b(n3624) );
	inv_2 U1308 ( .x(n1910), .a(N2007) );
	inv_2 U1309 ( .x(n1913), .a(N1941) );
	nand2i_2 U131 ( .x(n4010), .a(n694), .b(n891) );
	nand2i_2 U1310 ( .x(n1400), .a(n1913), .b(n3662) );
	nor2i_3 U1311 ( .x(n1396), .a(n1397), .b(n1055) );
	aoi211_1 U1312 ( .x(n3119), .a(N1643), .b(n809), .c(n1395), .d(n1393) );
	inv_2 U1313 ( .x(n1911), .a(N1742) );
	nand2i_2 U1314 ( .x(n3120), .a(n1911), .b(___cell__39620_net145150) );
	and4i_3 U1315 ( .x(n1399), .a(n1396), .b(n3120), .c(n3121), .d(n3119) );
	aoi22_1 U1316 ( .x(n2796), .a(n2797), .b(n2022), .c(n513), .d(n2024) );
	nand2i_2 U1317 ( .x(n2800), .a(n702), .b(n570) );
	nand2i_2 U1318 ( .x(n2794), .a(n1824), .b(n2837) );
	inv_2 U1319 ( .x(n1824), .a(N327) );
	nand2_4 U132 ( .x(n2184), .a(n3354), .b(n1558) );
	ao22_3 U1320 ( .x(n2788), .a(n2902), .b(n649), .c(n2863), .d(n650) );
	nor2i_2 U1321 ( .x(n1266), .a(n1267), .b(n1268) );
	inv_5 U1322 ( .x(n3368), .a(n3365) );
	or3i_2 U1323 ( .x(n1265), .a(n2768), .b(n2767), .c(n1260) );
	oai22_1 U1324 ( .x(n2767), .a(___cell__39620_net143710), .b(n1828), .c(___cell__39620_net143660),
		.d(n1827) );
	inv_2 U1325 ( .x(n1828), .a(N1751) );
	inv_2 U1326 ( .x(n1827), .a(N1718) );
	nor2_1 U1327 ( .x(n1260), .a(n947), .b(n1261) );
	inv_2 U1328 ( .x(n1261), .a(N1883) );
	inv_2 U1329 ( .x(n1833), .a(N2016) );
	ao22_4 U133 ( .x(n1999), .a(n627), .b(n3584), .c(n3448), .d(n659) );
	nand2i_2 U1330 ( .x(n1264), .a(n1833), .b(n3624) );
	inv_2 U1331 ( .x(n1829), .a(N1950) );
	nand2i_2 U1332 ( .x(n1263), .a(n1829), .b(n3662) );
	inv_8 U1333 ( .x(n2774), .a(n3856) );
	inv_2 U1334 ( .x(n1832), .a(N1983) );
	nand2i_2 U1335 ( .x(n2777), .a(n1832), .b(___cell__39620_net145508) );
	inv_2 U1336 ( .x(n1831), .a(N1850) );
	nand2i_2 U1337 ( .x(n2776), .a(n1831), .b(n4000) );
	inv_2 U1338 ( .x(n1830), .a(N1817) );
	nand2i_2 U1339 ( .x(n2775), .a(n1830), .b(n1987) );
	nand2i_2 U134 ( .x(n3701), .a(n4009), .b(n3196) );
	nand2i_2 U1340 ( .x(n3046), .a(n1588), .b(n3001) );
	aoi221_2 U1341 ( .x(n3039), .a(___cell__39620_net143864), .b(n3040), .c(n649),
		.d(n3041), .e(n3042) );
	aoi22_1 U1342 ( .x(n3050), .a(n2024), .b(n3012), .c(n1267), .d(n3051) );
	aoi21_1 U1343 ( .x(n3049), .a(n2022), .b(n3008), .c(n1359) );
	inv_2 U1344 ( .x(n3055), .a(n3964) );
	aoi21_1 U1345 ( .x(n3052), .a(n502), .b(n3054), .c(n3055) );
	nand2i_2 U1346 ( .x(n3047), .a(n1884), .b(n977) );
	inv_2 U1347 ( .x(n1884), .a(N354) );
	inv_2 U1348 ( .x(n1889), .a(N1844) );
	nand2i_2 U1349 ( .x(n3031), .a(n1889), .b(n4000) );
	aoi21_1 U135 ( .x(n2186), .a(n1249), .b(n2187), .c(n1121) );
	aoi22_1 U1350 ( .x(n3028), .a(N1811), .b(n1987), .c(n662), .d(n1339) );
	inv_2 U1351 ( .x(n1890), .a(N1977) );
	nand2i_2 U1352 ( .x(n3030), .a(n1890), .b(___cell__39620_net145508) );
	nand2i_2 U1353 ( .x(n1354), .a(n1885), .b(n3624) );
	inv_2 U1354 ( .x(n1885), .a(N2010) );
	inv_2 U1355 ( .x(n1888), .a(N1944) );
	nand2i_2 U1356 ( .x(n1353), .a(n1888), .b(n3999) );
	nor2i_1 U1357 ( .x(n1351), .a(N1745), .b(___cell__39620_net143710) );
	nand4i_1 U1358 ( .x(n3024), .a(n1350), .b(n3025), .c(n3026), .d(n3027) );
	nand4i_3 U1359 ( .x(n2989), .a(n1323), .b(n3937), .c(n3936), .d(n3935) );
	oai22_1 U136 ( .x(n2230), .a(n1570), .b(n1715), .c(n512), .d(n1713) );
	inv_2 U1360 ( .x(n3079), .a(n3973) );
	nand2i_2 U1361 ( .x(n3086), .a(n1892), .b(n977) );
	inv_2 U1362 ( .x(n1892), .a(N353) );
	ao21_3 U1363 ( .x(n3083), .a(n2022), .b(n3051), .c(n1374) );
	aoi21_1 U1364 ( .x(n3067), .a(n1197), .b(n1380), .c(n1364) );
	inv_2 U1365 ( .x(n1898), .a(N1976) );
	nand2i_2 U1366 ( .x(n3066), .a(n1898), .b(___cell__39620_net145508) );
	inv_2 U1367 ( .x(n1897), .a(N1810) );
	nand2i_2 U1368 ( .x(n3065), .a(n1897), .b(n1987) );
	nand2i_2 U1369 ( .x(n1367), .a(n1893), .b(n3624) );
	aoi21_1 U137 ( .x(n2231), .a(n1256), .b(n2130), .c(n2230) );
	inv_2 U1370 ( .x(n1893), .a(N2009) );
	inv_2 U1371 ( .x(n1896), .a(N1943) );
	nand2i_2 U1372 ( .x(n1366), .a(n1896), .b(n3662) );
	nor2i_1 U1373 ( .x(n1363), .a(N1744), .b(___cell__39620_net143710) );
	inv_2 U1374 ( .x(n1894), .a(N1645) );
	oai211_1 U1375 ( .x(n3062), .a(___cell__39620_net143872), .b(n1894), .c(n3061),
		.d(n3063) );
	inv_2 U1376 ( .x(___cell__39620_net144347), .a(___cell__39620_net144343) );
	aoi211_1 U1377 ( .x(n1365), .a(n1318), .b(n594), .c(n3062), .d(n1363) );
	inv_5 U1378 ( .x(n2011), .a(n2054) );
	nand2i_2 U1379 ( .x(n3163), .a(n1917), .b(n2837) );
	inv_8 U138 ( .x(n1686), .a(n1684) );
	inv_2 U1380 ( .x(n1917), .a(N317) );
	nand2i_2 U1381 ( .x(n3162), .a(n1588), .b(n2014) );
	aoai211_1 U1382 ( .x(n3158), .a(n1217), .b(n3159), .c(n1572), .d(n3155) );
	aoi21_1 U1383 ( .x(n3173), .a(n3174), .b(n1085), .c(n1415) );
	aoi221_1 U1384 ( .x(n3167), .a(n2022), .b(n3168), .c(n1267), .d(n2023),
		.e(n1414) );
	nand2i_2 U1385 ( .x(n3164), .a(n1916), .b(n1064) );
	nand2i_2 U1386 ( .x(n3983), .a(n1918), .b(n977) );
	inv_2 U1387 ( .x(n1918), .a(N350) );
	aoi21_1 U1388 ( .x(n3153), .a(n1197), .b(n1054), .c(n1409) );
	inv_2 U1389 ( .x(n1922), .a(N1807) );
	nand2_2 U139 ( .x(n1712), .a(n1686), .b(___cell__39620_net144517) );
	nand2i_2 U1390 ( .x(n3154), .a(n1922), .b(n1987) );
	aoi22_1 U1391 ( .x(n3150), .a(n662), .b(n4141), .c(n1095), .d(n1992) );
	nand3_1 U1392 ( .x(n1413), .a(n3150), .b(n3154), .c(n3153) );
	nand2i_2 U1393 ( .x(n1412), .a(n1919), .b(n3624) );
	inv_2 U1394 ( .x(n1919), .a(N2006) );
	inv_2 U1395 ( .x(n1921), .a(N1940) );
	nand2i_2 U1396 ( .x(n1411), .a(n1921), .b(n3999) );
	ao21_3 U1397 ( .x(n3149), .a(n1318), .b(n1988), .c(n1408) );
	inv_2 U1398 ( .x(n1923), .a(N1973) );
	nand2i_2 U1399 ( .x(n3152), .a(n1923), .b(___cell__39620_net145508) );
	oai22_1 U140 ( .x(n2176), .a(n1584), .b(n1712), .c(n2177), .d(n1711) );
	aoi211_1 U1400 ( .x(n3148), .a(N1642), .b(n809), .c(n1407), .d(n1405) );
	inv_2 U1401 ( .x(n1920), .a(N1873) );
	nand2i_2 U1402 ( .x(n3151), .a(n1920), .b(n3998) );
	nand2i_2 U1403 ( .x(n2717), .a(n1658), .b(n3830) );
	nand2_2 U1404 ( .x(n2716), .a(n1085), .b(n3835) );
	nand2i_2 U1405 ( .x(n2704), .a(n1808), .b(n2837) );
	inv_2 U1406 ( .x(n1808), .a(N329) );
	inv_2 U1407 ( .x(n2699), .a(n3849) );
	nand2i_2 U1408 ( .x(n2702), .a(n1186), .b(n2574) );
	nor2i_3 U1409 ( .x(n2703), .a(n2709), .b(n2706) );
	aoi21_1 U141 ( .x(n2113), .a(n2070), .b(n583), .c(n1982) );
	nand2i_2 U1410 ( .x(n2685), .a(n1616), .b(n3839) );
	nand2i_2 U1411 ( .x(n2687), .a(n1815), .b(___cell__39620_net145508) );
	inv_2 U1412 ( .x(n1815), .a(N1985) );
	nand2i_2 U1413 ( .x(n2688), .a(n1814), .b(n735) );
	inv_2 U1414 ( .x(n1814), .a(N1852) );
	nand4i_1 U1415 ( .x(n2678), .a(n1240), .b(n2679), .c(n2680), .d(n2681) );
	inv_2 U1416 ( .x(n1810), .a(N2018) );
	nand2i_2 U1417 ( .x(n2684), .a(n1810), .b(n3624) );
	inv_2 U1418 ( .x(n1812), .a(N1885) );
	nand2i_2 U1419 ( .x(n2683), .a(n1812), .b(n944) );
	nand2_2 U142 ( .x(n2114), .a(n2115), .b(n2113) );
	and4i_3 U1420 ( .x(n1246), .a(n2678), .b(n2682), .c(n2683), .d(n2684) );
	inv_2 U1421 ( .x(n1813), .a(N1952) );
	nand2i_2 U1422 ( .x(n1245), .a(n1813), .b(n3999) );
	inv_2 U1423 ( .x(n1243), .a(N1819) );
	nor2_1 U1424 ( .x(n1242), .a(n1077), .b(n1243) );
	inv_2 U1425 ( .x(___cell__39620_net143785), .a(___cell__39620_net144350) );
	nand2i_2 U1426 ( .x(n2199), .a(n1588), .b(n2089) );
	aoi22_1 U1427 ( .x(n2196), .a(n650), .b(n2197), .c(n1221), .d(n2090) );
	aoi222_2 U1428 ( .x(n2191), .a(n649), .b(n2192), .c(n2193), .d(n2194),
		.e(n2139), .f(n2195) );
	nand4_1 U1429 ( .x(n2198), .a(n2191), .b(n2188), .c(n2196), .d(n2199) );
	inv_2 U143 ( .x(n664), .a(___cell__39620_net144326) );
	nand2i_2 U1430 ( .x(n2201), .a(n1703), .b(n977) );
	inv_2 U1431 ( .x(n1703), .a(N345) );
	and4i_3 U1432 ( .x(n2200), .a(n2209), .b(n2207), .c(n2202), .d(n2208) );
	nand2i_2 U1433 ( .x(n2207), .a(n670), .b(n3693) );
	inv_2 U1434 ( .x(n1705), .a(N1637) );
	nand2i_2 U1435 ( .x(n2170), .a(n1705), .b(n809) );
	inv_2 U1436 ( .x(n1706), .a(N1703) );
	nand2i_2 U1437 ( .x(n2169), .a(n1706), .b(___cell__39620_net145190) );
	aoi22_1 U1438 ( .x(n2166), .a(n1318), .b(n2167), .c(n1197), .d(n2168) );
	nand4_1 U1439 ( .x(n1129), .a(n2166), .b(n2164), .c(n2169), .d(n2170) );
	aoi21_1 U144 ( .x(n2069), .a(n2070), .b(n636), .c(n1982) );
	nand2i_2 U1440 ( .x(n1128), .a(n1704), .b(n3624) );
	inv_2 U1441 ( .x(n1704), .a(N2001) );
	inv_2 U1442 ( .x(n1708), .a(N1935) );
	nand2i_2 U1443 ( .x(n1127), .a(n1708), .b(n3662) );
	inv_2 U1444 ( .x(n1709), .a(N1968) );
	nand2i_2 U1445 ( .x(n2175), .a(n1709), .b(___cell__39620_net145508) );
	aoi22_1 U1446 ( .x(n2174), .a(N1802), .b(n1987), .c(N1835), .d(n4000) );
	inv_2 U1447 ( .x(n1707), .a(N1736) );
	nand2i_2 U1448 ( .x(n2173), .a(n1707), .b(___cell__39620_net145150) );
	aoi221_1 U1449 ( .x(n2862), .a(n1191), .b(n2863), .c(n1221), .d(n743),
		.e(n1297) );
	nand2i_0 U145 ( .x(n3706), .a(n1561), .b(n2070) );
	aoi22_1 U1450 ( .x(n2855), .a(n887), .b(n2856), .c(n502), .d(n2857) );
	inv_2 U1451 ( .x(n2861), .a(n1498) );
	inv_2 U1452 ( .x(n2860), .a(n1497) );
	aoi222_1 U1453 ( .x(n2858), .a(n649), .b(n2859), .c(n2193), .d(n2860),
		.e(n2139), .f(n2861) );
	aoi221_1 U1454 ( .x(n2871), .a(n2872), .b(n2022), .c(n842), .d(n2024),
		.e(n2869) );
	nand2i_2 U1456 ( .x(n2867), .a(n1844), .b(n2837) );
	inv_2 U1457 ( .x(n1844), .a(N326) );
	inv_2 U1458 ( .x(n1850), .a(N1982) );
	nand2i_2 U1459 ( .x(n2848), .a(n1850), .b(___cell__39620_net145508) );
	nand2i_2 U146 ( .x(n3707), .a(___cell__39620_net144317), .b(n1361) );
	aoi21_1 U1460 ( .x(n2845), .a(n1095), .b(n2846), .c(n1291) );
	inv_2 U1461 ( .x(n1848), .a(N1882) );
	nand2i_2 U1462 ( .x(n2847), .a(n1848), .b(n3998) );
	nand4_1 U1463 ( .x(n1296), .a(n2842), .b(n2847), .c(n2845), .d(n2848) );
	aoi221_1 U1464 ( .x(n1295), .a(n1197), .b(n2849), .c(N1849), .d(n735),
		.e(n1293) );
	inv_2 U1465 ( .x(n1849), .a(N1949) );
	nand2i_2 U1466 ( .x(n1294), .a(n1849), .b(n3999) );
	nand2i_2 U1467 ( .x(n2243), .a(n1574), .b(n2192) );
	aoi22_1 U1468 ( .x(n2241), .a(n1191), .b(n2197), .c(n1221), .d(n2089) );
	aoi221_1 U1469 ( .x(n2234), .a(n2211), .b(n2235), .c(n2212), .d(n750),
		.e(n1142) );
	inv_14 U147 ( .x(n940), .a(n938) );
	inv_2 U1470 ( .x(n2240), .a(n1468) );
	inv_2 U1471 ( .x(n2239), .a(n1467) );
	aoi222_1 U1472 ( .x(n2237), .a(n649), .b(n2238), .c(n2193), .d(n2239),
		.e(n2139), .f(n2240) );
	nand4_1 U1473 ( .x(n2242), .a(n2237), .b(n2234), .c(n2241), .d(n2243) );
	inv_2 U1474 ( .x(n1717), .a(N344) );
	nand2i_2 U1475 ( .x(n2244), .a(n1717), .b(n977) );
	inv_2 U1476 ( .x(n1718), .a(N1636) );
	nand2i_2 U1477 ( .x(n2221), .a(n1718), .b(n809) );
	aoi22_2 U1478 ( .x(n2219), .a(n1197), .b(n2165), .c(n662), .d(n2167) );
	nand2i_2 U1479 ( .x(n1140), .a(n1725), .b(n3624) );
	inv_5 U148 ( .x(n783), .a(Imm[0]) );
	inv_2 U1480 ( .x(n1725), .a(N2000) );
	inv_2 U1481 ( .x(n1721), .a(N1934) );
	nand2i_2 U1482 ( .x(n1139), .a(n1721), .b(n3999) );
	and4i_1 U1483 ( .x(n1138), .a(n2222), .b(n2223), .c(n2224), .d(n2225) );
	nand2i_2 U1484 ( .x(n2223), .a(n1722), .b(n1987) );
	inv_2 U1485 ( .x(n1722), .a(N1801) );
	nand2i_2 U1486 ( .x(n2224), .a(n1723), .b(n735) );
	inv_2 U1487 ( .x(n1723), .a(N1834) );
	nand2i_2 U1488 ( .x(n2225), .a(n1724), .b(___cell__39620_net145508) );
	inv_2 U1489 ( .x(n1724), .a(N1967) );
	nand2i_2 U149 ( .x(n3298), .a(n1579), .b(n928) );
	oai22_1 U1490 ( .x(n2222), .a(n947), .b(n1720), .c(___cell__39620_net143710),
		.d(n1719) );
	inv_2 U1491 ( .x(n1720), .a(N1867) );
	inv_2 U1492 ( .x(n1719), .a(N1735) );
	nand2i_2 U1493 ( .x(n2909), .a(n1852), .b(n2837) );
	inv_2 U1494 ( .x(n1852), .a(N325) );
	inv_5 U1495 ( .x(n633), .a(n632) );
	and3i_2 U1496 ( .x(n2905), .a(n2908), .b(n2906), .c(n2907) );
	nand2i_2 U1499 ( .x(n2904), .a(n1574), .b(n2859) );
	inv_10 U150 ( .x(n863), .a(n862) );
	and4i_2 U1500 ( .x(n2883), .a(n1307), .b(n2884), .c(n2885), .d(n2886) );
	nand2i_2 U1501 ( .x(n2884), .a(n1856), .b(___cell__39620_net145508) );
	inv_2 U1502 ( .x(n1856), .a(N1981) );
	oai22_2 U1503 ( .x(n2880), .a(n2774), .b(n1182), .c(n865), .d(n1055) );
	nor2i_3 U1504 ( .x(n1304), .a(N1749), .b(___cell__39620_net143710) );
	inv_2 U1505 ( .x(n1319), .a(n2846) );
	aoi221_1 U1506 ( .x(n2882), .a(n1197), .b(n2846), .c(N1848), .d(n4000),
		.e(n1305) );
	nor2i_1 U1507 ( .x(n1309), .a(N2014), .b(n1169) );
	and4i_4 U1508 ( .x(n2308), .a(___cell__39620_net143784), .b(n2311), .c(n2309),
		.d(n2310) );
	nand2_2 U151 ( .x(n3789), .a(n3478), .b(___cell__39620_net144331) );
	nand2i_4 U1510 ( .x(n3745), .a(n1736), .b(n944) );
	inv_2 U1511 ( .x(n821), .a(n1161) );
	inv_2 U1512 ( .x(n2328), .a(n3749) );
	aoi21_1 U1513 ( .x(n2327), .a(n1191), .b(n1728), .c(n2328) );
	nand2i_2 U1514 ( .x(n2331), .a(n703), .b(___cell__39620_net147270) );
	nand4i_1 U1515 ( .x(n2329), .a(n2330), .b(n2331), .c(n2332), .d(n2327) );
	aoi22_1 U1516 ( .x(n2317), .a(n535), .b(n2318), .c(___cell__39620_net143864),
		.d(n2319) );
	aoi21_1 U1517 ( .x(n2323), .a(___cell__39620_net143722), .b(n2324), .c(n2320) );
	nand2i_2 U1518 ( .x(n2326), .a(n2300), .b(n3741) );
	inv_2 U1519 ( .x(___cell__39620_net145472), .a(___cell__39620_net144555) );
	aoi22_1 U152 ( .x(n706), .a(n710), .b(n709), .c(n708), .d(n707) );
	aoi22_1 U1520 ( .x(___cell__39620_net145470), .a(___cell__39620_net145450),
		.b(n798), .c(___cell__39620_net145451), .d(___cell__39620_net145472) );
	inv_2 U1521 ( .x(n3776), .a(n1477) );
	nand2_2 U1522 ( .x(n2441), .a(n2193), .b(n3776) );
	nand2i_2 U1523 ( .x(n2440), .a(n1478), .b(n2139) );
	oai211_2 U1524 ( .x(n2438), .a(n2439), .b(n1658), .c(n2440), .d(n2441) );
	nand3i_2 U1525 ( .x(n2442), .a(n2443), .b(n2444), .c(n2445) );
	aoi21_1 U1526 ( .x(n2444), .a(n1221), .b(n2402), .c(n1190) );
	aoi22_1 U1527 ( .x(n2454), .a(reg_out_B[28]), .b(n1064), .c(Imm[28]), .d(___cell__39620_net145617) );
	aoi21_1 U1528 ( .x(n2453), .a(n2457), .b(___cell__39620_net143864), .c(n1192) );
	nand2i_2 U1529 ( .x(n2452), .a(___cell__39620_net144406), .b(n2499) );
	nand2_5 U153 ( .x(n615), .a(N1662), .b(n616) );
	aoi22_1 U1530 ( .x(n2451), .a(n2022), .b(n2455), .c(n2024), .d(n2456) );
	nand2i_2 U1531 ( .x(n2420), .a(n588), .b(n663) );
	inv_2 U1532 ( .x(n1757), .a(N1726) );
	nand2i_2 U1533 ( .x(n2419), .a(n1757), .b(___cell__39620_net145190) );
	nor2i_1 U1534 ( .x(n1188), .a(N1759), .b(___cell__39620_net143710) );
	nand4i_1 U1535 ( .x(n2418), .a(n1188), .b(n2419), .c(n2420), .d(n2421) );
	inv_2 U1536 ( .x(n1755), .a(N2024) );
	nand2i_2 U1537 ( .x(n2417), .a(n1755), .b(n3624) );
	inv_2 U1538 ( .x(n1756), .a(N1660) );
	nand2i_2 U1539 ( .x(n2416), .a(n1756), .b(n809) );
	inv_2 U154 ( .x(n3269), .a(n1472) );
	nand2i_2 U1540 ( .x(n2415), .a(n2412), .b(___cell__39620_net145285) );
	nand2i_2 U1541 ( .x(n2414), .a(n1182), .b(n3727) );
	nand4_1 U1542 ( .x(n2413), .a(n2414), .b(n2415), .c(n2416), .d(n2417) );
	inv_2 U1543 ( .x(n1758), .a(N1958) );
	nand2i_4 U1544 ( .x(n2427), .a(n1758), .b(n3662) );
	inv_2 U1545 ( .x(n1759), .a(N1825) );
	aoi22_1 U1547 ( .x(n2057), .a(n1267), .b(n2059), .c(n2024), .d(n2027) );
	nand2i_1 U1548 ( .x(n2052), .a(n1566), .b(n2090) );
	inv_5 U1549 ( .x(n3614), .a(n3613) );
	exnor2_1 U155 ( .x(n1472), .a(reg_out_A[30]), .b(reg_out_B[30]) );
	oai211_1 U1550 ( .x(n2051), .a(n2012), .b(n1574), .c(n2052), .d(n2049) );
	inv_2 U1551 ( .x(n1670), .a(N1971) );
	nand2i_2 U1552 ( .x(n2042), .a(n1670), .b(___cell__39620_net145508) );
	aoi21_2 U1553 ( .x(n2039), .a(n662), .b(n1054), .c(n1076) );
	inv_2 U1554 ( .x(n1669), .a(N1838) );
	nand2i_2 U1555 ( .x(n2041), .a(n1669), .b(n735) );
	aoi22_1 U1556 ( .x(n2040), .a(n1197), .b(n1993), .c(n1095), .d(n2043) );
	inv_2 U1557 ( .x(n1666), .a(N2004) );
	nand2i_2 U1558 ( .x(n2038), .a(n1666), .b(n3624) );
	aoi211_1 U1559 ( .x(n2035), .a(N1640), .b(n809), .c(n1075), .d(n1073) );
	exnor2_1 U156 ( .x(n1471), .a(reg_out_A[30]), .b(Imm[30]) );
	inv_2 U1560 ( .x(n1667), .a(N1871) );
	nand2i_2 U1561 ( .x(n2037), .a(n1667), .b(n944) );
	aoi22_1 U1562 ( .x(n2036), .a(N1739), .b(___cell__39620_net145150), .c(n1318),
		.d(n1992) );
	nand4_1 U1563 ( .x(n1080), .a(n2036), .b(n2037), .c(n2035), .d(n2038) );
	inv_2 U1564 ( .x(n1668), .a(N1938) );
	nand2i_2 U1565 ( .x(n1079), .a(n1668), .b(n3999) );
	inv_2 U1566 ( .x(n2400), .a(n578) );
	aoi221_1 U1567 ( .x(n2395), .a(n649), .b(n2399), .c(n650), .d(n2400), .e(n2396) );
	nand2i_2 U1568 ( .x(n2394), .a(n702), .b(n2324) );
	inv_2 U1569 ( .x(n2393), .a(n2319) );
	nand2i_2 U157 ( .x(n3775), .a(n1752), .b(n1063) );
	inv_2 U1571 ( .x(n3740), .a(n2402) );
	nand4i_1 U1572 ( .x(n2403), .a(n2405), .b(n2407), .c(n2408), .d(n2409) );
	aoi211_1 U1573 ( .x(n2401), .a(n1191), .b(n2402), .c(n2403), .d(n1185) );
	inv_7 U1574 ( .x(n3724), .a(n3723) );
	nand2i_2 U1576 ( .x(n2404), .a(n784), .b(n3765) );
	oai21_2 U1577 ( .x(n2391), .a(n816), .b(n3720), .c(n2372) );
	inv_2 U1578 ( .x(n3767), .a(n3766) );
	nand2i_2 U1579 ( .x(n2390), .a(n3767), .b(n1217) );
	inv_2 U158 ( .x(n2185), .a(n1715) );
	aoi22_1 U1580 ( .x(n2389), .a(n539), .b(n2390), .c(___cell__39620_net143722),
		.d(n2391) );
	nand4_1 U1581 ( .x(n2377), .a(n2378), .b(n2379), .c(n2380), .d(n2381) );
	nand2i_2 U1582 ( .x(n2378), .a(n1055), .b(n3727) );
	nand2i_2 U1583 ( .x(n2379), .a(n2376), .b(___cell__39620_net147791) );
	nand2i_2 U1584 ( .x(n2381), .a(n1750), .b(n3624) );
	inv_2 U1585 ( .x(n1750), .a(N2025) );
	aoi221_1 U1587 ( .x(n2383), .a(n1197), .b(n2384), .c(N1992), .d(___cell__39620_net145508),
		.e(n1181) );
	aoi21_1 U1588 ( .x(n791), .a(n535), .b(___cell__39620_net145444), .c(n782) );
	inv_7 U1589 ( .x(n3720), .a(n3719) );
	inv_2 U1590 ( .x(n792), .a(___cell__39620_net147270) );
	inv_2 U1591 ( .x(n798), .a(n794) );
	nand2_2 U1592 ( .x(___cell__39620_net145428), .a(n2288), .b(n2289) );
	inv_2 U1593 ( .x(n1727), .a(N1961) );
	inv_2 U1594 ( .x(___cell__39620_net144355), .a(___cell__39620_net143653) );
	inv_5 U1595 ( .x(___cell__39620_net143872), .a(n809) );
	inv_4 U1596 ( .x(n1726), .a(N2027) );
	oai21_1 U1597 ( .x(n2293), .a(n1153), .b(n1658), .c(n2294) );
	inv_2 U1598 ( .x(n678), .a(n1662) );
	nand3_3 U1599 ( .x(n1087), .a(n678), .b(n1663), .c(n701) );
	oai22_1 U160 ( .x(n2428), .a(n1529), .b(n1715), .c(n2429), .d(n1713) );
	nand4i_1 U1600 ( .x(n3988), .a(n1424), .b(n3190), .c(n3987), .d(n3192) );
	nor2i_1 U1601 ( .x(n1424), .a(N1997), .b(n1169) );
	nand2i_2 U1602 ( .x(n3987), .a(___cell__39620_net144343), .b(n3245) );
	inv_2 U1603 ( .x(n1426), .a(n1517) );
	nor2i_1 U1604 ( .x(n1425), .a(n1426), .b(n690) );
	ao21_2 U1605 ( .x(n3207), .a(n2024), .b(n2826), .c(n1425) );
	nand2i_2 U1606 ( .x(n3209), .a(n1518), .b(n2139) );
	nand2i_3 U1607 ( .x(n3206), .a(n1626), .b(n2827) );
	aoai211_1 U1608 ( .x(n3205), .a(n917), .b(n530), .c(n1064), .d(n816) );
	nand2i_0 U1609 ( .x(n3180), .a(___cell__39620_net144175), .b(n1545) );
	inv_5 U161 ( .x(n938), .a(reg_out_A[2]) );
	nand2i_2 U1610 ( .x(n3989), .a(n1924), .b(n2837) );
	inv_2 U1611 ( .x(n1924), .a(N308) );
	inv_5 U1612 ( .x(n1437), .a(n3219) );
	inv_5 U1613 ( .x(n3216), .a(n1733) );
	oai211_1 U1614 ( .x(n3215), .a(n3216), .b(n1657), .c(n3217), .d(n3218) );
	inv_5 U1615 ( .x(n941), .a(reg_out_A[0]) );
	aoi222_1 U1616 ( .x(n3212), .a(n502), .b(n3214), .c(n942), .d(___cell__39620_net145444),
		.e(N341), .f(n977) );
	inv_5 U1617 ( .x(n3611), .a(n3610) );
	inv_5 U1618 ( .x(n2012), .a(n2093) );
	nand2i_2 U1619 ( .x(n2016), .a(n1594), .b(n2837) );
	exnor2_1 U162 ( .x(n1475), .a(reg_out_A[29]), .b(Imm[29]) );
	inv_2 U1620 ( .x(n1594), .a(N316) );
	aoi21_1 U1622 ( .x(n2013), .a(n1221), .b(n2014), .c(n2007) );
	inv_2 U1623 ( .x(n3623), .a(n3622) );
	inv_5 U1624 ( .x(n3620), .a(n3619) );
	oai211_1 U1625 ( .x(n2007), .a(n1062), .b(n1532), .c(n2008), .d(n2009) );
	aoi22_1 U1626 ( .x(n2026), .a(n502), .b(n2027), .c(___cell__39620_net143722),
		.d(n2028) );
	inv_2 U1627 ( .x(n2025), .a(n720) );
	aoi22_1 U1628 ( .x(n2021), .a(n2022), .b(n2023), .c(n2024), .d(n2025) );
	nand3_1 U1629 ( .x(n2020), .a(n2021), .b(n2029), .c(n2026) );
	inv_2 U163 ( .x(n3266), .a(n1476) );
	nand2i_2 U1630 ( .x(n2019), .a(n1598), .b(n977) );
	inv_2 U1631 ( .x(n1598), .a(N349) );
	nand2i_2 U1633 ( .x(n2033), .a(n1658), .b(n3172) );
	inv_2 U1634 ( .x(n1615), .a(N1839) );
	nand2i_2 U1635 ( .x(n1991), .a(n1615), .b(n4000) );
	aoi22_1 U1636 ( .x(n1986), .a(N1806), .b(n1987), .c(n662), .d(n1988) );
	inv_2 U1637 ( .x(n1617), .a(N1972) );
	nand2i_2 U1638 ( .x(n1990), .a(n1617), .b(___cell__39620_net145508) );
	aoi22_1 U1639 ( .x(n1989), .a(n1197), .b(n1992), .c(n1095), .d(n1993) );
	nand2_5 U164 ( .x(n1089), .a(n713), .b(n927) );
	nand2i_2 U1640 ( .x(n1058), .a(n1599), .b(n3624) );
	inv_2 U1641 ( .x(n1599), .a(N2005) );
	inv_2 U1642 ( .x(n1613), .a(N1939) );
	nand2i_2 U1643 ( .x(n1057), .a(n1613), .b(n3662) );
	and4i_3 U1644 ( .x(n1056), .a(n1053), .b(n1984), .c(n1985), .d(n1983) );
	nand2i_2 U1645 ( .x(n1984), .a(n1600), .b(___cell__39620_net145150) );
	inv_2 U1646 ( .x(n1600), .a(N1740) );
	nand2i_2 U1647 ( .x(n1985), .a(n1601), .b(n3998) );
	inv_2 U1648 ( .x(n1601), .a(N1872) );
	aoi211_1 U1649 ( .x(n1983), .a(N1641), .b(n809), .c(n1052), .d(n1050) );
	nand2i_1 U165 ( .x(___cell__39620_net144555), .a(n498), .b(n1728) );
	aoi22_1 U1650 ( .x(n3011), .a(n502), .b(n3012), .c(___cell__39620_net143722),
		.d(n3013) );
	aoi21_1 U1651 ( .x(n3003), .a(n1191), .b(n3004), .c(___cell__39620_net143982) );
	aoi22_1 U1652 ( .x(n2999), .a(n649), .b(n3000), .c(n650), .d(n3001) );
	aoi21_1 U1653 ( .x(n3002), .a(n1221), .b(n2899), .c(n2996) );
	inv_2 U1654 ( .x(n1876), .a(N355) );
	nand2i_2 U1655 ( .x(n3006), .a(n1876), .b(n977) );
	nand2i_4 U1656 ( .x(n2987), .a(n1881), .b(n735) );
	aoi21_1 U1657 ( .x(n2985), .a(n662), .b(n1308), .c(n1340) );
	inv_4 U1658 ( .x(n1882), .a(N1978) );
	nand2i_4 U1659 ( .x(n2986), .a(n1882), .b(___cell__39620_net145508) );
	nand2i_2 U166 ( .x(n3761), .a(n1635), .b(___cell__39620_net145472) );
	nand2i_2 U1660 ( .x(n1344), .a(n1877), .b(n3624) );
	inv_2 U1661 ( .x(n1877), .a(N2011) );
	inv_2 U1662 ( .x(n1880), .a(N1945) );
	nand2i_2 U1663 ( .x(n1343), .a(n1880), .b(n3662) );
	inv_2 U1664 ( .x(n1879), .a(N1878) );
	inv_2 U1665 ( .x(n1878), .a(N1746) );
	nand2i_2 U1666 ( .x(n2983), .a(n1878), .b(___cell__39620_net145150) );
	aoi211_1 U1667 ( .x(n2982), .a(N1647), .b(n809), .c(n1337), .d(n1335) );
	inv_2 U1668 ( .x(n1868), .a(N356) );
	aoi21_1 U1669 ( .x(n2965), .a(n1191), .b(n2899), .c(n1327) );
	nand2i_2 U167 ( .x(___cell__39620_net147350), .a(n718), .b(n798) );
	nand2i_2 U1670 ( .x(n2970), .a(n1867), .b(n2837) );
	inv_2 U1671 ( .x(n1867), .a(N323) );
	nand2i_2 U1672 ( .x(n2963), .a(n1574), .b(n3004) );
	and3i_1 U1673 ( .x(n2962), .a(n2961), .b(n2963), .c(n2964) );
	inv_2 U1674 ( .x(n1871), .a(N1946) );
	nand2i_2 U1675 ( .x(n3938), .a(n1871), .b(n3662) );
	inv_2 U1676 ( .x(n1873), .a(N2012) );
	nand2i_2 U1677 ( .x(n3939), .a(n1873), .b(n3624) );
	nand4_1 U1678 ( .x(n2954), .a(n2955), .b(n2956), .c(n2957), .d(n2953) );
	nand4i_1 U1679 ( .x(n3940), .a(n2954), .b(n2950), .c(n3939), .d(n3938) );
	or2_1 U168 ( .x(n498), .a(reg_out_B[4]), .b(reg_out_B[3]) );
	nand4i_1 U1680 ( .x(n3912), .a(n2920), .b(n2918), .c(n3910), .d(n3911) );
	nand4_1 U1681 ( .x(n2920), .a(n2921), .b(n2922), .c(n2923), .d(n2924) );
	nand2i_2 U1682 ( .x(n3910), .a(n1863), .b(n3999) );
	inv_2 U1683 ( .x(n1863), .a(N1947) );
	nand2i_2 U1684 ( .x(n3911), .a(n1865), .b(n3624) );
	inv_2 U1685 ( .x(n1865), .a(N2013) );
	nand3i_1 U1686 ( .x(n2931), .a(n2932), .b(n2933), .c(n2934) );
	nand2i_2 U1687 ( .x(n2947), .a(n1857), .b(n2837) );
	inv_2 U1688 ( .x(n1857), .a(N324) );
	nand2i_2 U1689 ( .x(n2946), .a(n1858), .b(n977) );
	inv_5 U169 ( .x(___cell__39620_net144707), .a(Imm[24]) );
	inv_2 U1690 ( .x(n1858), .a(N357) );
	nand2i_2 U1691 ( .x(n2752), .a(n1817), .b(n2837) );
	inv_2 U1692 ( .x(n1817), .a(N328) );
	nor3i_2 U1693 ( .x(n2749), .a(n2747), .b(n2748), .c(n2745) );
	inv_2 U1694 ( .x(n1816), .a(n567) );
	ao22_3 U1695 ( .x(n2759), .a(n757), .b(n2803), .c(n3854), .d(n758) );
	nand2i_2 U1696 ( .x(n2761), .a(n4001), .b(n2714) );
	and3i_3 U1697 ( .x(n2750), .a(n2759), .b(n2760), .c(n2761) );
	nand4i_2 U1698 ( .x(n2724), .a(n2723), .b(n2725), .c(n2726), .d(n2727) );
	inv_2 U1699 ( .x(n1821), .a(N1884) );
	inv_5 U170 ( .x(n648), .a(Imm[29]) );
	nand2i_2 U1700 ( .x(n2736), .a(n1821), .b(n3997) );
	aoi21_1 U1701 ( .x(n2732), .a(n1197), .b(n2733), .c(n1253) );
	inv_2 U1702 ( .x(n1818), .a(N1653) );
	nand2i_2 U1703 ( .x(n2735), .a(n1818), .b(n809) );
	and4i_3 U1704 ( .x(n2734), .a(n2724), .b(n2735), .c(n2732), .d(n2736) );
	nand2i_4 U1705 ( .x(n2731), .a(n1822), .b(n3662) );
	inv_2 U1706 ( .x(n1823), .a(N1818) );
	nand2i_2 U1707 ( .x(n2730), .a(n1823), .b(n1987) );
	nand4i_1 U1708 ( .x(n2728), .a(n1251), .b(n2729), .c(n2730), .d(n2731) );
	nor2i_1 U1709 ( .x(n1252), .a(N2017), .b(n1169) );
	exnor2_1 U171 ( .x(n1470), .a(reg_out_A[31]), .b(n4144) );
	inv_2 U1710 ( .x(n2668), .a(n3835) );
	inv_5 U1711 ( .x(n3553), .a(n3552) );
	nand2i_2 U1712 ( .x(n2671), .a(n4030), .b(n3057) );
	nand4_1 U1713 ( .x(n2624), .a(n3825), .b(n3824), .c(n3823), .d(n3822) );
	aoi22_1 U1714 ( .x(n2660), .a(n829), .b(___cell__39620_net145617), .c(n2661),
		.d(n2024) );
	nand2_2 U1715 ( .x(n2663), .a(n2707), .b(n502) );
	nand4_1 U1716 ( .x(n2662), .a(n2663), .b(n2664), .c(n2660), .d(n2665) );
	buf_10 U1717 ( .x(n636), .a(reg_out_A[23]) );
	inv_2 U1718 ( .x(n3841), .a(n3840) );
	inv_2 U1719 ( .x(n2652), .a(n1488) );
	nor2i_1 U172 ( .x(n1149), .a(n1150), .b(n509) );
	inv_2 U1720 ( .x(n2651), .a(n1487) );
	aoi22_1 U1721 ( .x(n2650), .a(n2139), .b(n2651), .c(n2193), .d(n2652) );
	oai211_3 U1722 ( .x(n3837), .a(n747), .b(n1565), .c(n3836), .d(n2628) );
	inv_5 U1723 ( .x(n2655), .a(n3837) );
	oai211_1 U1724 ( .x(n2654), .a(n2655), .b(n1566), .c(n2650), .d(n2656) );
	nand2i_2 U1725 ( .x(n2659), .a(n1798), .b(n2837) );
	inv_2 U1726 ( .x(n1798), .a(N330) );
	nand2i_2 U1727 ( .x(n3842), .a(n1797), .b(n1064) );
	inv_2 U1728 ( .x(n2658), .a(n3842) );
	oai221_4 U1729 ( .x(n2574), .a(n3419), .b(n1070), .c(n1313), .d(n1565),
		.e(n1807) );
	nand2_1 U173 ( .x(n3401), .a(n1691), .b(n901) );
	aoi21_1 U1730 ( .x(n2657), .a(n1191), .b(n2574), .c(n2658) );
	inv_2 U1731 ( .x(n1800), .a(N2019) );
	nand2i_2 U1732 ( .x(n2642), .a(n1800), .b(n3624) );
	inv_2 U1733 ( .x(n1803), .a(N1886) );
	nand2i_2 U1734 ( .x(n2641), .a(n1803), .b(n3998) );
	inv_2 U1735 ( .x(n1802), .a(N1721) );
	nand2i_2 U1736 ( .x(n2640), .a(n1802), .b(___cell__39620_net145190) );
	and4i_1 U1737 ( .x(n1239), .a(n2636), .b(n2640), .c(n2641), .d(n2642) );
	nand2i_2 U1738 ( .x(n2647), .a(n1804), .b(n3999) );
	aoi211_1 U1739 ( .x(n2646), .a(n1197), .b(n2600), .c(n1237), .d(n1236) );
	nand2i_3 U174 ( .x(n3729), .a(n1564), .b(n3591) );
	nand2i_2 U1740 ( .x(n2627), .a(n1658), .b(n3812) );
	nand2_2 U1741 ( .x(n2626), .a(n1085), .b(n3816) );
	nand2i_2 U1742 ( .x(n2625), .a(n4031), .b(n3057) );
	nand4_1 U1743 ( .x(n2618), .a(n2625), .b(n2626), .c(n2623), .d(n2627) );
	inv_2 U1744 ( .x(n1791), .a(N364) );
	nand2i_2 U1745 ( .x(n2617), .a(n1791), .b(n977) );
	inv_5 U1746 ( .x(n2611), .a(n3422) );
	inv_2 U1747 ( .x(n1790), .a(N331) );
	nand2i_2 U1748 ( .x(n3827), .a(n1790), .b(n2837) );
	inv_2 U1749 ( .x(n2615), .a(n3827) );
	aoi22_1 U175 ( .x(n2269), .a(n1971), .b(n2270), .c(n1177), .d(n2271) );
	inv_2 U1750 ( .x(n2613), .a(n3828) );
	nor3i_2 U1751 ( .x(n2614), .a(n2612), .b(n2615), .c(n2610) );
	nand2_2 U1752 ( .x(n2621), .a(n2661), .b(n502) );
	and4i_3 U1753 ( .x(n1232), .a(n2598), .b(n2596), .c(n2592), .d(n2597) );
	nand2i_2 U1754 ( .x(n2596), .a(n1796), .b(___cell__39620_net145508) );
	inv_2 U1755 ( .x(n1796), .a(N1987) );
	and4i_3 U1756 ( .x(n2592), .a(n2589), .b(n2593), .c(n2594), .d(n2595) );
	nand2i_2 U1757 ( .x(n1231), .a(n1792), .b(n3624) );
	inv_2 U1758 ( .x(n1792), .a(N2020) );
	nand2i_2 U1759 ( .x(n2559), .a(n1788), .b(n3999) );
	inv_3 U176 ( .x(n3462), .a(n2265) );
	aoi221_1 U1760 ( .x(n2555), .a(n1318), .b(n2473), .c(n662), .d(n2423),
		.e(n1213) );
	nor2i_3 U1761 ( .x(n1215), .a(N1988), .b(___cell__39620_net143845) );
	nand4i_1 U1762 ( .x(n2558), .a(n1215), .b(n2555), .c(n2556), .d(n2559) );
	inv_2 U1763 ( .x(n1784), .a(N2021) );
	nand2i_2 U1764 ( .x(n2554), .a(n1784), .b(n3624) );
	inv_2 U1765 ( .x(n1787), .a(N1888) );
	nand2i_2 U1766 ( .x(n2553), .a(n1787), .b(n944) );
	inv_2 U1767 ( .x(n1786), .a(N1723) );
	nand2i_2 U1768 ( .x(n2552), .a(n1786), .b(___cell__39620_net145190) );
	inv_2 U1769 ( .x(n2550), .a(n3819) );
	nand2i_2 U177 ( .x(n2265), .a(n3492), .b(n3493) );
	and4i_1 U1770 ( .x(n2547), .a(n2550), .b(n2548), .c(n2549), .d(n2546) );
	nand4_1 U1771 ( .x(n2551), .a(n2547), .b(n2552), .c(n2553), .d(n2554) );
	nand2i_2 U1772 ( .x(n1454), .a(n1060), .b(n1591) );
	nand2i_2 U1773 ( .x(n2587), .a(n784), .b(n3812) );
	inv_2 U1774 ( .x(n2586), .a(n3816) );
	oai211_2 U1775 ( .x(n2579), .a(n2586), .b(___cell__39620_net144406), .c(n2580),
		.d(n2587) );
	aoi22_1 U1776 ( .x(n2573), .a(n649), .b(n2574), .c(n650), .d(n2532) );
	aoi21_1 U1777 ( .x(n2567), .a(n2544), .b(n2568), .c(n1216) );
	nor2i_3 U1778 ( .x(n1223), .a(n1204), .b(n1224) );
	nand2i_2 U1779 ( .x(n2585), .a(n4032), .b(n3057) );
	aoi22_1 U178 ( .x(n2264), .a(n2079), .b(n2265), .c(n2266), .d(n608) );
	nand2i_2 U1780 ( .x(n2542), .a(n4001), .b(n3782) );
	nand2i_2 U1781 ( .x(n2541), .a(n4033), .b(n3057) );
	inv_2 U1782 ( .x(n2540), .a(n3785) );
	oai211_1 U1783 ( .x(n2538), .a(n2540), .b(n702), .c(n2541), .d(n2542) );
	nand2i_2 U1784 ( .x(n2537), .a(n1772), .b(n2837) );
	inv_2 U1785 ( .x(n1710), .a(n1447) );
	aoi22_1 U1786 ( .x(n2536), .a(reg_out_B[26]), .b(n1064), .c(Imm[26]), .d(___cell__39620_net145617) );
	nor2i_3 U1787 ( .x(n1210), .a(___cell__39620_net143722), .b(n1211) );
	inv_2 U1788 ( .x(n1591), .a(n1590) );
	nand2i_2 U1789 ( .x(n1595), .a(n1534), .b(n1591) );
	inv_2 U1790 ( .x(n1597), .a(n1595) );
	inv_2 U1791 ( .x(n3805), .a(n3804) );
	inv_2 U1792 ( .x(n3807), .a(n3806) );
	aoai211_1 U1793 ( .x(n2529), .a(n502), .b(n2568), .c(n3807), .d(n1451) );
	inv_4 U1794 ( .x(n3809), .a(n3808) );
	inv_2 U1795 ( .x(n2524), .a(n2489) );
	oai211_1 U1796 ( .x(n2523), .a(n2524), .b(n1580), .c(n2525), .d(n2526) );
	nand4i_3 U1797 ( .x(n2527), .a(n2523), .b(n2528), .c(n2529), .d(n2530) );
	inv_2 U1798 ( .x(n3420), .a(n2673) );
	aoi22_1 U1799 ( .x(n2531), .a(n539), .b(n2490), .c(n649), .d(n2532) );
	nand2i_2 U180 ( .x(n2263), .a(n1625), .b(n2302) );
	inv_2 U1800 ( .x(n3423), .a(n3739) );
	nand2i_2 U1801 ( .x(n2534), .a(n1574), .b(n3422) );
	inv_8 U1802 ( .x(n3418), .a(n2763) );
	aoi22_1 U1803 ( .x(n2533), .a(n1221), .b(n2399), .c(n1191), .d(n2492) );
	inv_8 U1804 ( .x(n1520), .a(n1519) );
	nand3_1 U1805 ( .x(n1184), .a(n1520), .b(n810), .c(n1612) );
	nor2i_1 U1806 ( .x(n1209), .a(N1956), .b(n1184) );
	inv_2 U1807 ( .x(n1774), .a(N2022) );
	nand2i_2 U1808 ( .x(n2511), .a(n1774), .b(n3624) );
	inv_2 U1809 ( .x(n1777), .a(N1889) );
	nand2i_2 U181 ( .x(n3734), .a(n1564), .b(n3594) );
	nand2i_2 U1810 ( .x(n2510), .a(n1777), .b(n3998) );
	inv_4 U1811 ( .x(n1776), .a(N1724) );
	nand2i_3 U1812 ( .x(n2509), .a(n1776), .b(___cell__39620_net145190) );
	inv_2 U1813 ( .x(n2507), .a(n3803) );
	nand2i_2 U1814 ( .x(n2515), .a(n1616), .b(n2473) );
	inv_2 U1815 ( .x(n1779), .a(N1989) );
	nand2i_2 U1816 ( .x(n2517), .a(n1780), .b(n4000) );
	nor2i_1 U1817 ( .x(___cell__39620_net144312), .a(___cell__39620_net144166),
		.b(n805) );
	aoi211_1 U1818 ( .x(n1005), .a(n977), .b(N343), .c(n2364), .d(n2354) );
	oai211_1 U1819 ( .x(n4052), .a(n1004), .b(___cell__39620_net147731), .c(n1005),
		.d(n1006) );
	nor2i_3 U182 ( .x(n1151), .a(n1147), .b(n1152) );
	aoi221_1 U1820 ( .x(n953), .a(N309), .b(n2837), .c(N342), .d(n977), .e(n2834) );
	ao21_2 U1821 ( .x(n4055), .a(___cell__39620_net143326), .b(n999), .c(n1000) );
	inv_2 U1822 ( .x(n1899), .a(N319) );
	nand2i_2 U1823 ( .x(n968), .a(n1899), .b(n2837) );
	inv_2 U1824 ( .x(n1674), .a(N314) );
	nand2i_2 U1825 ( .x(n959), .a(n1674), .b(n2837) );
	and4i_3 U1826 ( .x(n989), .a(n2497), .b(n2495), .c(n2493), .d(n2496) );
	inv_2 U1827 ( .x(n1762), .a(N367) );
	nand2i_2 U1828 ( .x(n988), .a(n1762), .b(n977) );
	nand2i_2 U1829 ( .x(n1456), .a(n4018), .b(n3057) );
	oai21_1 U183 ( .x(n2259), .a(n1529), .b(n1281), .c(n2260) );
	and4i_1 U1830 ( .x(n1036), .a(n3129), .b(n3132), .c(n3133), .d(n3134) );
	inv_2 U1831 ( .x(n1825), .a(N360) );
	nand2i_2 U1832 ( .x(n1022), .a(n1825), .b(n977) );
	and4i_3 U1833 ( .x(n1021), .a(n2795), .b(n2793), .c(n2792), .d(n2794) );
	and4i_2 U1834 ( .x(n1020), .a(n1265), .b(n1262), .c(n1263), .d(n1264) );
	inv_2 U1836 ( .x(n1883), .a(N321) );
	nand2i_2 U1837 ( .x(n971), .a(n1883), .b(n2837) );
	inv_2 U1838 ( .x(n1891), .a(N320) );
	nand2i_2 U1839 ( .x(n1032), .a(n1891), .b(n2837) );
	nor2_0 U184 ( .x(n1938), .a(IR_function_field[4]), .b(IR_function_field[1]) );
	and4i_1 U1840 ( .x(n965), .a(n3160), .b(n3161), .c(n3162), .d(n3163) );
	inv_2 U1841 ( .x(n1809), .a(N362) );
	nand2i_2 U1842 ( .x(n1019), .a(n1809), .b(n977) );
	and4i_3 U1843 ( .x(n1018), .a(n2705), .b(n2703), .c(n2700), .d(n2704) );
	and4i_2 U1844 ( .x(n1017), .a(n1247), .b(n1244), .c(n1245), .d(n1246) );
	inv_2 U1845 ( .x(n1702), .a(N312) );
	nand2i_2 U1846 ( .x(n956), .a(n1702), .b(n2837) );
	and4i_2 U1847 ( .x(n954), .a(n1129), .b(n1126), .c(n1127), .d(n1128) );
	inv_2 U1848 ( .x(n1845), .a(N359) );
	nand2i_2 U1849 ( .x(n1025), .a(n1845), .b(n977) );
	inv_4 U185 ( .x(n3861), .a(n1834) );
	nor3i_2 U1850 ( .x(n1024), .a(n2867), .b(n2868), .c(n2865) );
	and3i_2 U1851 ( .x(n1023), .a(n1296), .b(n1294), .c(n1295) );
	inv_2 U1852 ( .x(n1716), .a(N311) );
	nand2i_2 U1853 ( .x(n1003), .a(n1716), .b(n2837) );
	oai211_1 U1854 ( .x(n4053), .a(n1001), .b(___cell__39620_net143287), .c(n1002),
		.d(n1003) );
	inv_2 U1855 ( .x(n1853), .a(N358) );
	nand2i_2 U1856 ( .x(n3891), .a(n1853), .b(n977) );
	inv_2 U1857 ( .x(n976), .a(n3891) );
	nand4_1 U1858 ( .x(n975), .a(n2905), .b(n2896), .c(n2903), .d(n2909) );
	inv_2 U1860 ( .x(n859), .a(n2329) );
	inv_2 U1861 ( .x(n1753), .a(N335) );
	nand2i_2 U1862 ( .x(n1007), .a(n1753), .b(n2837) );
	inv_2 U1863 ( .x(n1754), .a(N368) );
	nand2i_4 U1864 ( .x(n1009), .a(n1754), .b(n977) );
	inv_2 U1866 ( .x(n1665), .a(N315) );
	nand2i_2 U1867 ( .x(n997), .a(n1665), .b(n2837) );
	nor3i_1 U1868 ( .x(n996), .a(n1079), .b(n1080), .c(n1081) );
	oai31_2 U1869 ( .x(n993), .a(n2387), .b(n2377), .c(n2382), .d(___cell__39620_net147732) );
	oaoi211_1 U187 ( .x(n1416), .a(n1417), .b(n1418), .c(n665), .d(___cell__39620_net144062) );
	nand2i_2 U1870 ( .x(n991), .a(n1748), .b(n2837) );
	inv_2 U1871 ( .x(n1748), .a(N336) );
	nand3i_1 U1872 ( .x(n1942), .a(IR_opcode_field[0]), .b(n1533), .c(___cell__39620_net143655) );
	inv_2 U1873 ( .x(n3211), .a(n3989) );
	nand3i_1 U1874 ( .x(n948), .a(n3211), .b(n3212), .c(n3213) );
	inv_2 U1875 ( .x(n1875), .a(N322) );
	nand2i_2 U1876 ( .x(n1030), .a(n1875), .b(n2837) );
	nand2i_2 U1877 ( .x(n972), .a(___cell__39620_net143287), .b(n3940) );
	and4i_4 U1878 ( .x(n1026), .a(n2937), .b(n2940), .c(n2946), .d(n2947) );
	nand2i_2 U1879 ( .x(n1027), .a(___cell__39620_net147731), .b(n3912) );
	inv_2 U188 ( .x(n1421), .a(N1864) );
	or3i_2 U1880 ( .x(n978), .a(n2734), .b(n1252), .c(n2728) );
	inv_8 U1881 ( .x(n807), .a(n806) );
	inv_2 U1882 ( .x(n1799), .a(N363) );
	nand2i_2 U1883 ( .x(n981), .a(n1799), .b(n977) );
	oai21_1 U1884 ( .x(n986), .a(n2551), .b(n2558), .c(___cell__39620_net143326) );
	inv_2 U1885 ( .x(n1783), .a(N365) );
	nand2i_2 U1886 ( .x(n985), .a(n1783), .b(n977) );
	inv_2 U1887 ( .x(n1782), .a(N332) );
	nand2i_2 U1888 ( .x(n984), .a(n1782), .b(n2837) );
	nand2i_2 U1889 ( .x(n1013), .a(n1773), .b(n977) );
	nor2_1 U189 ( .x(n1420), .a(n947), .b(n1421) );
	inv_2 U1890 ( .x(n1773), .a(N366) );
	inv_2 U1891 ( .x(n1533), .a(n733) );
	aoi21_1 U1892 ( .x(n4117), .a(n3997), .b(n945), .c(___cell__6067_net21981) );
	nor2i_1 U1893 ( .x(N3297), .a(n4144), .b(n4116) );
	inv_2 U1894 ( .x(n1530), .a(IR_function_field[0]) );
	inv_5 U1895 ( .x(n744), .a(Imm[22]) );
	inv_2 U1896 ( .x(n1781), .a(reg_out_B[25]) );
	inv_2 U1897 ( .x(n1671), .a(n4146) );
	inv_2 U1899 ( .x(n1797), .a(reg_out_B[23]) );
	inv_2 U190 ( .x(n3558), .a(n3664) );
	inv_2 U1900 ( .x(n1523), .a(IR_function_field[2]) );
	inv_0 U1901 ( .x(n1664), .a(reg_out_B[8]) );
	inv_5 U1902 ( .x(n830), .a(Imm[23]) );
	inv_2 U1903 ( .x(n1752), .a(reg_out_B[28]) );
	inv_2 U1905 ( .x(N144), .a(Imm[31]) );
	inv_2 U1906 ( .x(N70), .a(reg_out_B[31]) );
	inv_8 U1907 ( .x(n653), .a(reg_out_B[12]) );
	or2_2 U1908 ( .x(n496), .a(reg_out_B[0]), .b(IR_function_field[0]) );
	or2_2 U1909 ( .x(n497), .a(IR_opcode_field[1]), .b(net152465) );
	nand2_2 U191 ( .x(n3559), .a(n665), .b(n3630) );
	aoi21_6 U1910 ( .x(n499), .a(n2890), .b(n1602), .c(n3532) );
	aoi21_4 U1911 ( .x(n500), .a(n1685), .b(n541), .c(n3558) );
	and2_3 U1912 ( .x(n501), .a(n549), .b(n548) );
	and2_8 U1913 ( .x(n502), .a(n619), .b(n1444) );
	inv_16 U1914 ( .x(n650), .a(n1574) );
	oa21_2 U1915 ( .x(n503), .a(net149120), .b(n517), .c(n4140) );
	inv_2 U1916 ( .x(n805), .a(n810) );
	and2_6 U1917 ( .x(n810), .a(n803), .b(IR_opcode_field[3]) );
	and2_8 U1918 ( .x(n504), .a(n726), .b(n725) );
	oaoi211_4 U1919 ( .x(n578), .a(n3585), .b(n575), .c(n576), .d(n577) );
	nand2i_2 U192 ( .x(n1418), .a(n1676), .b(___cell__39620_net144330) );
	inv_16 U1920 ( .x(n855), .a(reg_out_B[4]) );
	inv_2 U1921 ( .x(n675), .a(IR_opcode_field[1]) );
	or2_4 U1922 ( .x(n1524), .a(IR_function_field[1]), .b(IR_function_field[0]) );
	oa22_4 U1923 ( .x(n510), .a(n1580), .b(n1651), .c(n1578), .d(n890) );
	inv_2 U1924 ( .x(n1584), .a(n634) );
	buf_12 U1925 ( .x(n583), .a(reg_out_A[22]) );
	inv_2 U1926 ( .x(n3532), .a(n3758) );
	nand2i_2 U1927 ( .x(n3758), .a(n1655), .b(n811) );
	inv_2 U1928 ( .x(n671), .a(n891) );
	inv_12 U1929 ( .x(n748), .a(reg_out_A[20]) );
	nand2i_2 U193 ( .x(n3716), .a(n748), .b(n2070) );
	mux2_4 U1930 ( .x(n513), .d0(n3379), .sl(n729), .d1(n3374) );
	inv_5 U1931 ( .x(n3335), .a(n2133) );
	nand2i_2 U1932 ( .x(n3699), .a(n1693), .b(n977) );
	inv_14 U1933 ( .x(n834), .a(n833) );
	and2_1 U1934 ( .x(n514), .a(n675), .b(net152465) );
	aoi222_1 U1935 ( .x(n515), .a(n1267), .b(n3008), .c(n2022), .d(n3009),
		.e(n2024), .f(n3010) );
	or2_6 U1936 ( .x(n1043), .a(n637), .b(Imm[3]) );
	inv_2 U1937 ( .x(n1333), .a(n4005) );
	nand2i_8 U1938 ( .x(___cell__39620_net144170), .a(IR_opcode_field[0]),
		.b(n1520) );
	ao22_3 U1939 ( .x(n518), .a(n1095), .b(n2988), .c(n1197), .d(n2989) );
	nand2_2 U194 ( .x(n1837), .a(n2268), .b(n910) );
	ao21_4 U1940 ( .x(n519), .a(n1238), .b(n1239), .c(___cell__39620_net143287) );
	mux2i_1 U1941 ( .x(n2581), .d0(n3444), .sl(net149120), .d1(n3788) );
	inv_16 U1942 ( .x(n943), .a(n941) );
	oa22_4 U1943 ( .x(n520), .a(n1644), .b(n889), .c(n1646), .d(n1651) );
	ao22_6 U1944 ( .x(n521), .a(n858), .b(n3584), .c(n2184), .d(n857) );
	inv_2 U1945 ( .x(n3307), .a(n761) );
	inv_14 U1946 ( .x(n862), .a(reg_out_A[17]) );
	oai22_5 U1947 ( .x(n3019), .a(n1529), .b(n880), .c(n822), .d(n1657) );
	inv_7 U1948 ( .x(n3357), .a(n3019) );
	inv_0 U1949 ( .x(n523), .a(n930) );
	nand2_2 U195 ( .x(n3279), .a(n3554), .b(n3555) );
	inv_2 U1950 ( .x(n524), .a(n523) );
	oai22_1 U1951 ( .x(n525), .a(n880), .b(n1648), .c(n822), .d(n1647) );
	inv_14 U1952 ( .x(n880), .a(n1643) );
	inv_10 U1953 ( .x(n3366), .a(n3369) );
	oai22_6 U1954 ( .x(n3369), .a(n1580), .b(n1629), .c(n748), .d(n881) );
	nand4_1 U1955 ( .x(n2865), .a(n2858), .b(n2866), .c(n2855), .d(n2862) );
	aoi22_2 U1956 ( .x(n3098), .a(n1256), .b(n1997), .c(n1249), .d(n3036) );
	aoi22_2 U1957 ( .x(n3035), .a(n1714), .b(n1997), .c(n1256), .d(n3036) );
	nand2i_2 U1958 ( .x(n3918), .a(n4009), .b(n1997) );
	inv_2 U1959 ( .x(n1767), .a(N1890) );
	nand2_2 U196 ( .x(n3339), .a(n1691), .b(n749) );
	inv_2 U1960 ( .x(n526), .a(n3357) );
	inv_1 U1961 ( .x(n527), .a(n799) );
	aoi22_3 U1962 ( .x(n2925), .a(n1714), .b(n2851), .c(n1256), .d(n2852) );
	inv_5 U1963 ( .x(n538), .a(n1580) );
	inv_0 U1964 ( .x(n1874), .a(reg_out_B[15]) );
	exnor2_1 U1965 ( .x(n1505), .a(reg_out_B[15]), .b(n608) );
	nand2i_2 U1966 ( .x(n1956), .a(reg_out_B[15]), .b(n1955) );
	inv_0 U1967 ( .x(n1789), .a(reg_out_B[24]) );
	exnor2_1 U1968 ( .x(n1485), .a(n541), .b(reg_out_B[24]) );
	inv_8 U197 ( .x(n1691), .a(n1688) );
	and4i_2 U1970 ( .x(n1035), .a(n3138), .b(n3135), .c(n3136), .d(n3137) );
	and4i_3 U1971 ( .x(n1034), .a(n1402), .b(n1399), .c(n1400), .d(n1401) );
	inv_14 U1972 ( .x(n689), .a(n688) );
	aoi22_4 U1973 ( .x(n528), .a(reg_out_A[29]), .b(n529), .c(reg_out_A[21]),
		.d(n883) );
	inv_5 U1974 ( .x(n3302), .a(n528) );
	inv_12 U1975 ( .x(n530), .a(n646) );
	and2_8 U1976 ( .x(n531), .a(n532), .b(___cell__39620_net144317) );
	inv_6 U1977 ( .x(n532), .a(n1603) );
	inv_12 U1979 ( .x(n533), .a(n1587) );
	nand2i_2 U198 ( .x(n3690), .a(n1546), .b(n1968) );
	oai21_3 U1980 ( .x(n3992), .a(n1433), .b(n1944), .c(n810) );
	inv_16 U1981 ( .x(n536), .a(n1546) );
	aoi221_1 U1982 ( .x(n2569), .a(n2543), .b(n2570), .c(n538), .d(n2490),
		.e(n2571) );
	oai21_1 U1983 ( .x(n2449), .a(n1732), .b(n2410), .c(n538) );
	nand2_0 U1984 ( .x(n2412), .a(Imm[28]), .b(n538) );
	nand2i_2 U1985 ( .x(n1711), .a(___cell__39620_net144317), .b(___cell__39620_net144517) );
	nand2i_2 U1986 ( .x(n1682), .a(___cell__39620_net144317), .b(n1683) );
	nand2i_2 U1987 ( .x(n3694), .a(___cell__39620_net144317), .b(n1349) );
	nand2i_2 U1988 ( .x(n3717), .a(___cell__39620_net144317), .b(n1042) );
	inv_2 U1989 ( .x(n534), .a(___cell__39620_net144317) );
	inv_4 U199 ( .x(n935), .a(reg_out_A[6]) );
	inv_2 U1991 ( .x(n535), .a(___cell__39620_net144257) );
	inv_2 U1992 ( .x(___cell__39620_net144257), .a(reg_out_A[30]) );
	inv_5 U1993 ( .x(n1546), .a(reg_out_B[3]) );
	inv_2 U1994 ( .x(n537), .a(n1587) );
	inv_8 U1995 ( .x(n1580), .a(reg_out_A[28]) );
	inv_5 U1996 ( .x(n539), .a(n1564) );
	inv_5 U1997 ( .x(n1564), .a(reg_out_A[29]) );
	inv_10 U1998 ( .x(n3433), .a(n3602) );
	nand4i_2 U1999 ( .x(n2387), .a(n1183), .b(n2385), .c(n2383), .d(n2388) );
	nand2i_4 U200 ( .x(n3340), .a(n1649), .b(n883) );
	mx4_4 U2000 ( .x(n2382), .d0(N1727), .sl0(___cell__39620_net145190), .d1(n556),
		.sl1(n663), .d2(N1892), .sl2(n3998), .d3(N1760), .sl3(n562) );
	nor2i_1 U2001 ( .x(n1278), .a(n1177), .b(n1279) );
	inv_2 U2002 ( .x(n1279), .a(n3318) );
	inv_16 U2003 ( .x(n590), .a(n1219) );
	inv_5 U2004 ( .x(n540), .a(n1573) );
	inv_5 U2005 ( .x(n541), .a(n1578) );
	inv_2 U2006 ( .x(n543), .a(reset) );
	inv_2 U2007 ( .x(n542), .a(reset) );
	inv_2 U2008 ( .x(n4017), .a(reset) );
	aoi221_3 U2009 ( .x(n2313), .a(N1761), .b(___cell__39620_net145150), .c(N1728),
		.d(___cell__39620_net145190), .e(n613) );
	aoai211_1 U201 ( .x(n3179), .a(n2066), .b(n902), .c(n2067), .d(n504) );
	nand2_8 U2010 ( .x(n825), .a(n1630), .b(n1546) );
	oai211_1 U2011 ( .x(n544), .a(n3460), .b(n719), .c(n3858), .d(n2782) );
	nand2i_6 U2012 ( .x(n3858), .a(___cell__39620_net144062), .b(n2520) );
	oai211_3 U2013 ( .x(n2802), .a(n3460), .b(n719), .c(n3858), .d(n2782) );
	inv_10 U2014 ( .x(n1630), .a(n1556) );
	and3i_3 U2015 ( .x(n2017), .a(n2030), .b(n2033), .c(n2034) );
	oai211_4 U2016 ( .x(n2030), .a(n868), .b(n702), .c(n2031), .d(n2032) );
	aoi22_1 U2017 ( .x(n2906), .a(___cell__39620_net143722), .b(n2910), .c(___cell__39620_net143864),
		.d(n2911) );
	inv_2 U2018 ( .x(n546), .a(n545) );
	inv_14 U2019 ( .x(n889), .a(n888) );
	inv_2 U202 ( .x(n2160), .a(n3350) );
	nand2_2 U2020 ( .x(n779), .a(___cell__39620_net144029), .b(n780) );
	inv_10 U2021 ( .x(___cell__39620_net144029), .a(Imm[12]) );
	or3i_5 U2023 ( .x(n774), .a(n775), .b(Imm[7]), .c(Imm[30]) );
	ao22_6 U2024 ( .x(n3085), .a(n764), .b(n3112), .c(n3054), .d(n765) );
	mux2i_3 U2025 ( .x(n842), .d0(n856), .sl(n848), .d1(n3368) );
	aoi21_1 U2026 ( .x(n2232), .a(n1249), .b(n2233), .c(n1134) );
	nand2_1 U2027 ( .x(n3692), .a(n1256), .b(n2233) );
	nand2_1 U2028 ( .x(n3668), .a(n1714), .b(n2233) );
	buf_3 U2029 ( .x(n547), .a(n584) );
	inv_5 U203 ( .x(n1175), .a(n823) );
	and2_3 U2030 ( .x(n584), .a(n585), .b(n644) );
	nand4_1 U2031 ( .x(n4075), .a(n1014), .b(n1012), .c(n1013), .d(n1011) );
	inv_2 U2032 ( .x(n548), .a(n1577) );
	inv_5 U2033 ( .x(n1577), .a(n893) );
	inv_2 U2034 ( .x(n549), .a(n1603) );
	inv_5 U2035 ( .x(n1569), .a(n910) );
	and4i_5 U2036 ( .x(n1551), .a(n1960), .b(n1958), .c(n600), .d(n601) );
	inv_2 U2037 ( .x(n600), .a(n4139) );
	oai22_5 U2039 ( .x(n2520), .a(n1586), .b(n836), .c(n3391), .d(n4125) );
	nor2_1 U204 ( .x(n897), .a(n899), .b(n898) );
	oai211_3 U2040 ( .x(n1423), .a(n3506), .b(n1602), .c(n665), .d(n2812) );
	aoi21_3 U2041 ( .x(n2812), .a(n1147), .b(n1049), .c(n1834) );
	nand4_4 U2042 ( .x(n2938), .a(n3895), .b(n3894), .c(n3893), .d(n3892) );
	nand2i_6 U2043 ( .x(n3895), .a(n719), .b(n3069) );
	inv_5 U2044 ( .x(n551), .a(___cell__39620_net144781) );
	inv_5 U2045 ( .x(___cell__39620_net144781), .a(Imm[20]) );
	aoi21_3 U2046 ( .x(n2344), .a(n1147), .b(n1047), .c(n1738) );
	inv_16 U2047 ( .x(n3355), .a(n521) );
	inv_5 U2048 ( .x(n762), .a(n3416) );
	nor3_5 U2049 ( .x(n2940), .a(n2939), .b(n2941), .c(n2942) );
	oa22_3 U205 ( .x(n508), .a(n880), .b(n1648), .c(n822), .d(n1647) );
	nand2i_1 U2050 ( .x(n3871), .a(n4010), .b(n3483) );
	nand2i_3 U2051 ( .x(n3893), .a(n1623), .b(n3483) );
	aoi21_2 U2052 ( .x(n2747), .a(n1221), .b(n2609), .c(n2743) );
	aoi22_1 U2053 ( .x(n2653), .a(n1221), .b(n2532), .c(n650), .d(n2609) );
	aoi21_1 U2054 ( .x(n2698), .a(n1191), .b(n2609), .c(n2699) );
	nand3_0 U2055 ( .x(n552), .a(n810), .b(___cell__39620_net144166), .c(___cell__39620_net143655) );
	inv_2 U2056 ( .x(n3998), .a(n552) );
	inv_2 U2057 ( .x(___cell__39620_net144166), .a(IR_opcode_field[0]) );
	mux2i_3 U2058 ( .x(n3283), .d0(n1949), .sl(IR_function_field[2]), .d1(n1948) );
	inv_2 U206 ( .x(n3450), .a(n897) );
	nand4i_2 U2060 ( .x(n797), .a(___cell__39620_net147731), .b(n652), .c(n708),
		.d(N1994) );
	nand2i_4 U2061 ( .x(n2298), .a(n1596), .b(N371) );
	nand3_2 U2062 ( .x(n2910), .a(n3878), .b(n3877), .c(n2887) );
	aoi22_2 U2063 ( .x(n2887), .a(n1249), .b(n2888), .c(n1714), .d(n2690) );
	inv_6 U2064 ( .x(n769), .a(n704) );
	inv_14 U2065 ( .x(n839), .a(n569) );
	nand4_1 U2066 ( .x(n3108), .a(n3115), .b(n3114), .c(n3109), .d(n3111) );
	nand2i_8 U2067 ( .x(n3484), .a(n1584), .b(n928) );
	nand2_0 U2068 ( .x(n3644), .a(___cell__39620_net144330), .b(n533) );
	nand2_0 U2069 ( .x(n3652), .a(___cell__39620_net144330), .b(reg_out_A[30]) );
	nand2i_3 U207 ( .x(n3470), .a(n3471), .b(n3472) );
	oa21_6 U2070 ( .x(n553), .a(n3426), .b(n618), .c(n3572) );
	inv_10 U2071 ( .x(n2386), .a(n553) );
	aoi22_4 U2072 ( .x(n3070), .a(n1256), .b(n2994), .c(n1249), .d(n2995) );
	nand2_8 U2074 ( .x(n2798), .a(n2780), .b(n2778) );
	nor2i_1 U2075 ( .x(n554), .a(N370), .b(n1596) );
	nand2i_1 U2076 ( .x(n3825), .a(n1635), .b(n2433) );
	or2_5 U2077 ( .x(n992), .a(n1749), .b(n1596) );
	nand2i_8 U2078 ( .x(n1596), .a(___cell__39620_net144175), .b(n1597) );
	oai211_3 U2079 ( .x(n3219), .a(n840), .b(___cell__39620_net144345), .c(n3199),
		.d(n3200) );
	nand2i_3 U208 ( .x(n3321), .a(n3322), .b(n3323) );
	nand3i_1 U2080 ( .x(n1937), .a(n1521), .b(IR_function_field[3]), .c(n1938) );
	mux2i_1 U2081 ( .x(n3593), .d0(n1531), .sl(IR_function_field[3]), .d1(IR_function_field[4]) );
	or3i_3 U2082 ( .x(___cell__39620_net145426), .a(N1828), .b(___cell__39620_net147731),
		.c(n1077) );
	inv_2 U2084 ( .x(n556), .a(n555) );
	inv_2 U2085 ( .x(n557), .a(n627) );
	buf_16 U2086 ( .x(n838), .a(n937) );
	nand2i_2 U2087 ( .x(n3362), .a(n1583), .b(n928) );
	aoi22_1 U2088 ( .x(n3111), .a(n2024), .b(n3112), .c(n1267), .d(n3113) );
	inv_10 U209 ( .x(n871), .a(n3575) );
	nand2_5 U2090 ( .x(n1973), .a(n1040), .b(n1974) );
	nand2_5 U2091 ( .x(n3343), .a(n1040), .b(n3608) );
	nand2_5 U2092 ( .x(n3325), .a(n1040), .b(n3603) );
	nand2_5 U2093 ( .x(n3311), .a(n1040), .b(n3607) );
	nor2i_3 U2094 ( .x(n2213), .a(n1040), .b(n2214) );
	nor2i_3 U2095 ( .x(n2159), .a(n1040), .b(n2160) );
	oai21_1 U2096 ( .x(n3276), .a(n1577), .b(n1730), .c(n1040) );
	nand2i_8 U2097 ( .x(n1603), .a(___cell__39620_net144329), .b(___cell__39620_net144331) );
	inv_10 U2098 ( .x(n923), .a(n1603) );
	nand2i_4 U2099 ( .x(n3754), .a(n1602), .b(n3687) );
	oai22_1 U210 ( .x(n559), .a(n1569), .b(n871), .c(n4125), .d(n1283) );
	inv_16 U2100 ( .x(___cell__39620_net143997), .a(Imm[14]) );
	inv_2 U2101 ( .x(n3174), .a(n860) );
	oai22_2 U2102 ( .x(n3139), .a(___cell__39620_net144406), .b(n860), .c(n3140),
		.d(n621) );
	mux2i_3 U2103 ( .x(n860), .d0(n3410), .sl(n625), .d1(n850) );
	aoi21_2 U2104 ( .x(n2760), .a(n1085), .b(n2713), .c(n1254) );
	oai211_2 U2105 ( .x(n574), .a(n3656), .b(n1043), .c(n2675), .d(n3846) );
	oai211_3 U2106 ( .x(n4058), .a(n960), .b(___cell__39620_net143287), .c(n961),
		.d(n962) );
	and3i_3 U2107 ( .x(n1545), .a(n1541), .b(IR_function_field[0]), .c(n1448) );
	nand2i_2 U2108 ( .x(n3919), .a(n1634), .b(n3369) );
	nand2_6 U2109 ( .x(n1631), .a(n1630), .b(n1546) );
	ao211_4 U211 ( .x(n1042), .a(net151904), .b(n3481), .c(n3465), .d(n1982) );
	oai211_2 U2110 ( .x(n4063), .a(n969), .b(___cell__39620_net147731), .c(n970),
		.d(n971) );
	oai22_1 U2111 ( .x(n558), .a(n1569), .b(n871), .c(n4125), .d(n1283) );
	oai22_2 U2112 ( .x(n1995), .a(n1569), .b(n871), .c(n4125), .d(n1283) );
	nand2i_3 U2113 ( .x(n2715), .a(n4029), .b(n3057) );
	ao22_5 U2114 ( .x(n2187), .a(n3327), .b(n763), .c(n887), .d(n3584) );
	inv_2 U2115 ( .x(n1583), .a(n887) );
	exnor2_1 U2116 ( .x(n1498), .a(n887), .b(reg_out_B[19]) );
	nand2_2 U2117 ( .x(n1739), .a(n3573), .b(n887) );
	exnor2_1 U2118 ( .x(n1497), .a(n887), .b(n684) );
	nand2i_2 U2119 ( .x(n2421), .a(n947), .b(N1891) );
	nand2_2 U212 ( .x(n3480), .a(n665), .b(n3635) );
	and4i_4 U2120 ( .x(___cell__39620_net144322), .a(n778), .b(n560), .c(n561),
		.d(___cell__39620_net144707) );
	inv_2 U2121 ( .x(n560), .a(Imm[31]) );
	inv_2 U2122 ( .x(n561), .a(Imm[19]) );
	inv_2 U2123 ( .x(n562), .a(___cell__39620_net143710) );
	and3i_4 U2124 ( .x(___cell__39620_net144321), .a(n774), .b(n648), .c(n647) );
	inv_5 U2125 ( .x(n647), .a(Imm[28]) );
	nand2_1 U2126 ( .x(n2380), .a(n809), .b(N1661) );
	ao221_4 U2127 ( .x(n2209), .a(n2247), .b(n1267), .c(n3702), .d(n563), .e(n564) );
	inv_2 U2128 ( .x(n563), .a(n621) );
	inv_2 U2129 ( .x(n564), .a(n2210) );
	nand2_2 U213 ( .x(n3479), .a(n665), .b(n3653) );
	and4i_3 U2130 ( .x(n1016), .a(n2618), .b(n2616), .c(n2614), .d(n2617) );
	inv_10 U2131 ( .x(n884), .a(n623) );
	oai211_4 U2132 ( .x(n2753), .a(n670), .b(n2754), .c(n2755), .d(n2756) );
	nand2_2 U2133 ( .x(n2665), .a(n845), .b(n2022) );
	nand2_2 U2134 ( .x(n2622), .a(n845), .b(n1267) );
	mux2i_3 U2135 ( .x(n845), .d0(n846), .sl(net150405), .d1(n510) );
	oai22_6 U2136 ( .x(n2841), .a(n875), .b(n1182), .c(n2774), .d(n1055) );
	inv_5 U2138 ( .x(n831), .a(n830) );
	nor2_4 U2139 ( .x(___cell__39620_net143596), .a(n788), .b(n790) );
	nand2i_2 U214 ( .x(n3945), .a(n4010), .b(n3547) );
	buf_3 U2140 ( .x(n567), .a(n4139) );
	buf_3 U2141 ( .x(n566), .a(n4139) );
	nand4_3 U2142 ( .x(n3081), .a(n660), .b(n3074), .c(n3080), .d(n3077) );
	mux2i_2 U2143 ( .x(n3171), .d0(n3358), .sl(n816), .d1(n3313) );
	aoi22_3 U2144 ( .x(n1994), .a(n559), .b(n1683), .c(___cell__39620_net144517),
		.d(n1996) );
	inv_7 U2145 ( .x(n1067), .a(n1996) );
	inv_0 U2146 ( .x(n568), .a(n806) );
	nand2i_8 U2147 ( .x(n806), .a(___cell__39620_net144173), .b(n708) );
	nor2_1 U2148 ( .x(n1206), .a(n1087), .b(n4034) );
	inv_14 U2149 ( .x(n644), .a(n643) );
	nand2i_2 U215 ( .x(n3946), .a(n718), .b(n2927) );
	inv_4 U2150 ( .x(n643), .a(n934) );
	oai211_3 U2151 ( .x(n4076), .a(n987), .b(___cell__39620_net143287), .c(n988),
		.d(n989) );
	aoi21_1 U2152 ( .x(n2092), .a(n1191), .b(n2093), .c(n1105) );
	nand2_8 U2153 ( .x(n569), .a(n1555), .b(n855) );
	aoi21_2 U2154 ( .x(n2228), .a(n1391), .b(n558), .c(n2226) );
	aoi22_2 U2155 ( .x(n2126), .a(n1391), .b(n1996), .c(n1066), .d(n1995) );
	nand3_1 U2156 ( .x(n570), .a(n3853), .b(n3852), .c(n2737) );
	aoi21_2 U2157 ( .x(n2053), .a(n1191), .b(n2054), .c(n1083) );
	aoi21_1 U2158 ( .x(n2091), .a(n1221), .b(n2054), .c(n2085) );
	inv_10 U2159 ( .x(n1417), .a(reg_out_A[17]) );
	nand2i_2 U216 ( .x(n3947), .a(___cell__39620_net144062), .b(n2854) );
	inv_10 U2160 ( .x(n892), .a(reg_out_A[16]) );
	nand2i_1 U2161 ( .x(n3928), .a(n1632), .b(n3019) );
	ao221_5 U2162 ( .x(n2197), .a(n3602), .b(n572), .c(n3691), .d(n824), .e(n571) );
	inv_0 U2163 ( .x(n572), .a(n1562) );
	nand2i_4 U2164 ( .x(n3435), .a(n4004), .b(n1969) );
	nand2_4 U2165 ( .x(n1562), .a(n815), .b(reg_out_B[3]) );
	inv_5 U2166 ( .x(n3434), .a(n3691) );
	nand2i_6 U2167 ( .x(n3691), .a(n2111), .b(n3690) );
	nand2i_3 U2168 ( .x(n3602), .a(n3601), .b(n3598) );
	nand4_5 U2169 ( .x(n771), .a(n573), .b(___cell__39620_net144322), .c(n772),
		.d(___cell__39620_net144321) );
	and4_5 U2170 ( .x(n573), .a(n607), .b(n1980), .c(n1979), .d(n1978) );
	and3i_4 U2171 ( .x(n772), .a(n776), .b(___cell__39620_net145078), .c(___cell__39620_net145077) );
	nor2i_1 U2172 ( .x(n2003), .a(IR_function_field[5]), .b(IR_function_field[2]) );
	inv_2 U2173 ( .x(n1521), .a(IR_function_field[5]) );
	nand3i_3 U2174 ( .x(n2059), .a(n1065), .b(n3665), .c(n2044) );
	oai211_2 U2175 ( .x(n4071), .a(n1017), .b(___cell__39620_net147731), .c(n1018),
		.d(n1019) );
	inv_6 U2176 ( .x(n875), .a(n574) );
	inv_10 U2177 ( .x(n3460), .a(n3458) );
	inv_5 U2178 ( .x(n575), .a(n3742) );
	inv_2 U2179 ( .x(n576), .a(n1565) );
	nand2i_4 U218 ( .x(n3456), .a(n1584), .b(n3575) );
	inv_2 U2180 ( .x(n577), .a(n3571) );
	inv_16 U2181 ( .x(n3585), .a(n1558) );
	inv_5 U2183 ( .x(n579), .a(n2056) );
	aoi221_3 U2185 ( .x(n2424), .a(n1197), .b(n2386), .c(N1991), .d(___cell__39620_net145508),
		.e(n1189) );
	nand2i_4 U2186 ( .x(n2388), .a(n1751), .b(n4000) );
	nand2i_2 U2187 ( .x(n2408), .a(n4036), .b(n3057) );
	nor2i_3 U2188 ( .x(n1084), .a(n1085), .b(n878) );
	inv_2 U2189 ( .x(n2028), .a(n878) );
	inv_5 U219 ( .x(n1331), .a(n1976) );
	inv_10 U2190 ( .x(n3446), .a(n3445) );
	oai22_6 U2191 ( .x(n3445), .a(n889), .b(n1655), .c(n1651), .d(n1654) );
	mux2i_2 U2192 ( .x(n878), .d0(n3414), .sl(reg_out_B[1]), .d1(n3545) );
	nand4_1 U2193 ( .x(n3138), .a(n3145), .b(n3144), .c(n3146), .d(n3147) );
	aoi222_3 U2194 ( .x(n2278), .a(n1066), .b(n2279), .c(n2266), .d(n644),
		.e(n2079), .f(n2280) );
	inv_10 U2195 ( .x(n925), .a(n923) );
	aoi22_4 U2196 ( .x(n2602), .a(n1683), .b(n2303), .c(___cell__39620_net144517),
		.d(n2603) );
	and4i_3 U2198 ( .x(n580), .a(n581), .b(n3668), .c(n3667), .d(n3666) );
	inv_2 U2199 ( .x(n3669), .a(n580) );
	exnor2_1 U220 ( .x(n1506), .a(net151622), .b(n609) );
	and2_5 U2200 ( .x(n581), .a(n504), .b(n2130) );
	aoi22_4 U2201 ( .x(n2691), .a(n1683), .b(n2603), .c(___cell__39620_net144517),
		.d(n2520) );
	inv_10 U2202 ( .x(n903), .a(reg_out_A[9]) );
	nand2_2 U2203 ( .x(n3145), .a(n3118), .b(n1204) );
	mux2i_5 U2204 ( .x(n3118), .d0(n499), .sl(n694), .d1(n3531) );
	and4i_3 U2205 ( .x(n2842), .a(n2841), .b(n2843), .c(n2840), .d(n2844) );
	nand2i_2 U2206 ( .x(n2843), .a(n1847), .b(___cell__39620_net145150) );
	inv_6 U2207 ( .x(n3486), .a(n3654) );
	inv_6 U2208 ( .x(n1450), .a(n3862) );
	nand4i_2 U2209 ( .x(n3165), .a(n3166), .b(n3167), .c(n3173), .d(n3169) );
	inv_5 U221 ( .x(n3476), .a(n3577) );
	inv_8 U2210 ( .x(n751), .a(n3576) );
	mux2i_5 U2211 ( .x(n2064), .d0(n520), .sl(net150405), .d1(n3518) );
	nand2i_2 U2212 ( .x(n3198), .a(n1687), .b(n3448) );
	nand2_2 U2213 ( .x(n3448), .a(n3449), .b(n3450) );
	nand3_5 U2215 ( .x(___cell__39620_net143597), .a(___cell__39620_net143326),
		.b(n657), .c(N1894) );
	oai22_6 U2216 ( .x(n2994), .a(n1219), .b(n822), .c(n557), .d(n881) );
	nand2_5 U2217 ( .x(n3475), .a(n582), .b(n1981) );
	inv_7 U2218 ( .x(n582), .a(n3476) );
	aoi21_2 U2219 ( .x(n1981), .a(net151904), .b(___cell__39620_net144328),
		.c(n1982) );
	nand2i_2 U222 ( .x(n3914), .a(n1623), .b(n3303) );
	nand2i_2 U2220 ( .x(n3795), .a(n4010), .b(n2603) );
	nand2i_2 U2221 ( .x(n3770), .a(n1623), .b(n2603) );
	mux2_6 U2222 ( .x(n2708), .d0(n3443), .sl(net150620), .d1(n3533) );
	oai22_2 U2223 ( .x(n3443), .a(n1564), .b(n1651), .c(n1219), .d(n889) );
	oai22_5 U2224 ( .x(n3533), .a(n1587), .b(n1651), .c(n891), .d(n3485) );
	nand4_2 U2225 ( .x(n979), .a(n2750), .b(n2751), .c(n2749), .d(n2752) );
	inv_1 U2226 ( .x(n585), .a(n1603) );
	nand2i_3 U2228 ( .x(n3579), .a(n4008), .b(n2179) );
	nand2i_2 U2229 ( .x(n3678), .a(n719), .b(n2179) );
	nand2i_2 U223 ( .x(n3915), .a(n1625), .b(n3033) );
	aoi22_1 U2230 ( .x(n2336), .a(n1391), .b(n2179), .c(___cell__39620_net144517),
		.d(n2337) );
	aoi21_2 U2231 ( .x(n2178), .a(n1066), .b(n2179), .c(n2176) );
	inv_7 U2232 ( .x(n886), .a(reg_out_A[19]) );
	and4i_4 U2233 ( .x(n1100), .a(n1094), .b(n2073), .c(n2072), .d(n2071) );
	inv_0 U2235 ( .x(n587), .a(___cell__39620_net144029) );
	inv_2 U2236 ( .x(n588), .a(n587) );
	oa22_1 U2237 ( .x(n895), .a(n889), .b(n1656), .c(n1651), .d(n1657) );
	nand4_3 U2238 ( .x(n3746), .a(n2314), .b(n3745), .c(n2312), .d(n2308) );
	inv_10 U2239 ( .x(n1552), .a(n1547) );
	nand4i_4 U2240 ( .x(n1547), .a(n1548), .b(n1551), .c(n1550), .d(n1549) );
	oai21_5 U2241 ( .x(n2433), .a(n536), .b(n3310), .c(n3387) );
	inv_10 U2242 ( .x(n913), .a(reg_out_A[8]) );
	inv_1 U2243 ( .x(n851), .a(reg_out_A[7]) );
	oai22_6 U2244 ( .x(n2181), .a(n1583), .b(n871), .c(n4125), .d(n3324) );
	ao221_4 U2246 ( .x(n2619), .a(n592), .b(n3996), .c(n2022), .d(n2581), .e(n591) );
	inv_2 U2247 ( .x(n591), .a(n2620) );
	inv_0 U2248 ( .x(n592), .a(n670) );
	inv_6 U2249 ( .x(n2583), .a(n3996) );
	nand2i_2 U225 ( .x(n3916), .a(___cell__39620_net144062), .b(n4127) );
	mux2i_6 U2250 ( .x(n3996), .d0(n3385), .sl(n816), .d1(n3779) );
	or2_8 U2251 ( .x(n3576), .a(n4140), .b(n593) );
	inv_0 U2252 ( .x(n593), .a(net151904) );
	nand4i_5 U2254 ( .x(n594), .a(n1332), .b(n3954), .c(n3953), .d(n3952) );
	oai221_5 U2255 ( .x(n2512), .a(n1198), .b(n1055), .c(n553), .d(n1182),
		.e(n2513) );
	mux2i_3 U2256 ( .x(n2106), .d0(n520), .sl(n595), .d1(n3525) );
	inv_2 U2257 ( .x(n595), .a(net150620) );
	inv_5 U2258 ( .x(n3525), .a(n2235) );
	nand2i_2 U2259 ( .x(n2637), .a(n1182), .b(n565) );
	nand2i_2 U2260 ( .x(n2590), .a(n1055), .b(n3523) );
	nand2i_2 U2261 ( .x(n3819), .a(n1616), .b(n565) );
	nand2i_2 U2262 ( .x(n3803), .a(n1166), .b(n565) );
	oai21_5 U2263 ( .x(n1738), .a(n890), .b(n1654), .c(n1739) );
	aoi221_1 U2264 ( .x(n3190), .a(n662), .b(n2218), .c(n3181), .d(___cell__39620_net145285),
		.e(n3187) );
	aoi22_1 U2265 ( .x(n2813), .a(n2811), .b(___cell__39620_net145285), .c(n1318),
		.d(n2218) );
	aoi22_1 U2266 ( .x(n2345), .a(n2343), .b(___cell__39620_net147791), .c(n1197),
		.d(n2218) );
	aoi22_1 U2267 ( .x(n2217), .a(n2215), .b(___cell__39620_net145285), .c(n1095),
		.d(n2218) );
	inv_12 U2268 ( .x(n890), .a(n888) );
	nand2i_2 U227 ( .x(n3917), .a(___cell__39620_net144374), .b(n3034) );
	aoi211_1 U2270 ( .x(n1352), .a(n1318), .b(n2989), .c(n3024), .d(n1351) );
	aoi22_1 U2271 ( .x(n3064), .a(n662), .b(n2989), .c(n1095), .d(n4141) );
	nand2i_4 U2272 ( .x(n2956), .a(n1166), .b(n2989) );
	inv_2 U2273 ( .x(n597), .a(n1660) );
	inv_2 U2274 ( .x(n598), .a(n4001) );
	oai211_2 U2275 ( .x(n4068), .a(___cell__39620_net147731), .b(n1023), .c(n1024),
		.d(n1025) );
	buf_16 U2276 ( .x(n603), .a(n4015) );
	nand4_1 U2277 ( .x(n2149), .a(n2152), .b(n2151), .c(n2147), .d(n2150) );
	nand2_8 U2278 ( .x(n3582), .a(n604), .b(n2181) );
	inv_2 U2279 ( .x(n604), .a(___cell__39620_net144374) );
	oai22_5 U228 ( .x(n1997), .a(n1577), .b(n881), .c(n1578), .d(n822) );
	inv_12 U2280 ( .x(n3600), .a(n3599) );
	nand2i_4 U2281 ( .x(n606), .a(n738), .b(n531) );
	inv_5 U2282 ( .x(n738), .a(Imm[2]) );
	nand4_1 U2284 ( .x(n4072), .a(n519), .b(n980), .c(n981), .d(n982) );
	inv_5 U2285 ( .x(n607), .a(Imm[26]) );
	nand4_3 U2286 ( .x(n3539), .a(n3717), .b(n3716), .c(n2216), .d(n1419) );
	nand4i_2 U2287 ( .x(n1345), .a(n518), .b(n2986), .c(n2985), .d(n2987) );
	inv_5 U2289 ( .x(n879), .a(reg_out_B[1]) );
	nand2i_2 U229 ( .x(n3921), .a(n1635), .b(n3036) );
	and2_2 U2290 ( .x(n622), .a(reg_out_A[9]), .b(n923) );
	and4_5 U2291 ( .x(n1550), .a(n1962), .b(n656), .c(n1961), .d(n1760) );
	inv_5 U2292 ( .x(n1961), .a(n736) );
	inv_2 U2294 ( .x(n936), .a(n935) );
	or2_6 U2295 ( .x(n1519), .a(IR_opcode_field[4]), .b(IR_opcode_field[5]) );
	nor2_1 U2296 ( .x(n1086), .a(n679), .b(n4044) );
	nand2i_8 U2297 ( .x(n610), .a(n1605), .b(n1606) );
	nand4i_5 U2298 ( .x(n3723), .a(n2274), .b(n3721), .c(n2276), .d(n3722) );
	aoi221_1 U2299 ( .x(n2599), .a(n1095), .b(n2600), .c(n1197), .d(n2557),
		.e(n1228) );
	nand2i_2 U230 ( .x(n3927), .a(n1634), .b(n2888) );
	aoi21_1 U2300 ( .x(n1244), .a(n662), .b(n2557), .c(n1242) );
	aoi22_1 U2301 ( .x(n2556), .a(N1855), .b(n4000), .c(n1095), .d(n2557) );
	oai211_4 U2302 ( .x(n3856), .a(n3639), .b(n4005), .c(n2721), .d(n3855) );
	inv_0 U2303 ( .x(n611), .a(net156363) );
	inv_0 U2304 ( .x(n612), .a(n663) );
	or2_2 U2305 ( .x(n614), .a(n611), .b(n612) );
	inv_0 U2306 ( .x(n616), .a(n706) );
	aoi222_1 U2307 ( .x(n2840), .a(N1651), .b(n809), .c(n2839), .d(___cell__39620_net147791),
		.e(n663), .f(n534) );
	nor2i_3 U2308 ( .x(n617), .a(net149627), .b(n779) );
	inv_4 U2309 ( .x(n776), .a(n617) );
	nand2i_2 U231 ( .x(n3929), .a(n1635), .b(n3020) );
	inv_12 U2310 ( .x(net149627), .a(Imm[8]) );
	inv_2 U2311 ( .x(n618), .a(n1333) );
	inv_10 U2312 ( .x(n3426), .a(n3764) );
	and4i_5 U2313 ( .x(___cell__39620_net143595), .a(___cell__39620_net145427),
		.b(___cell__39620_net145418), .c(___cell__39620_net145426), .d(___cell__39620_net145425) );
	inv_10 U2314 ( .x(n3518), .a(n3516) );
	nand4i_5 U2315 ( .x(n2514), .a(n2512), .b(n2515), .c(n2516), .d(n2517) );
	and2_8 U2316 ( .x(n619), .a(n620), .b(n807) );
	inv_16 U2317 ( .x(___cell__39620_net144175), .a(n619) );
	nand2_8 U2318 ( .x(n621), .a(n619), .b(n1444) );
	inv_10 U2319 ( .x(n1444), .a(n1452) );
	inv_5 U232 ( .x(n3294), .a(n3291) );
	nand2_6 U2320 ( .x(___cell__6067_net21981), .a(n1037), .b(n1038) );
	nand2_2 U2321 ( .x(n3477), .a(n665), .b(n3652) );
	nand2_2 U2322 ( .x(n3478), .a(n665), .b(n3644) );
	inv_5 U2323 ( .x(n1038), .a(counter[0]) );
	oai22_1 U2324 ( .x(n2226), .a(n1570), .b(n1712), .c(n2227), .d(n1711) );
	oai22_6 U2325 ( .x(n3451), .a(n1570), .b(n836), .c(n4125), .d(n2227) );
	oai22_1 U2327 ( .x(n3233), .a(n1577), .b(n1091), .c(n500), .d(n1682) );
	and4i_4 U2328 ( .x(___cell__39620_net145418), .a(n769), .b(___cell__39620_net145421),
		.c(___cell__39620_net145419), .d(net150643) );
	oai221_4 U2329 ( .x(n623), .a(n3509), .b(n1607), .c(n624), .d(n3510), .e(n3511) );
	nand2i_2 U233 ( .x(n3922), .a(n1623), .b(n3291) );
	inv_2 U2330 ( .x(n624), .a(n671) );
	inv_4 U2331 ( .x(n3509), .a(n3646) );
	nand2i_1 U2332 ( .x(n3828), .a(n1789), .b(n1064) );
	nand2i_2 U2333 ( .x(n3826), .a(n1789), .b(n1063) );
	oai21_5 U2334 ( .x(___cell__39620_net147278), .a(n3724), .b(___cell__39620_net144345),
		.c(n2278) );
	oa22_5 U2335 ( .x(n2807), .a(n843), .b(n512), .c(n1175), .d(n1570) );
	and3i_3 U2336 ( .x(n1033), .a(n3081), .b(n3082), .c(n3086) );
	mux2i_5 U2337 ( .x(n3677), .d0(n3313), .sl(n625), .d1(n3314) );
	inv_2 U2338 ( .x(n625), .a(n739) );
	inv_0 U2339 ( .x(n626), .a(n4140) );
	nand2i_2 U234 ( .x(n3923), .a(n4010), .b(n2890) );
	nand2i_0 U2340 ( .x(n3136), .a(___cell__39620_net144655), .b(___cell__39620_net145617) );
	inv_0 U2341 ( .x(n627), .a(n1417) );
	inv_0 U2342 ( .x(n629), .a(n905) );
	oai211_1 U2344 ( .x(n4060), .a(n1034), .b(___cell__39620_net147731), .c(n1035),
		.d(n1036) );
	aoi21_1 U2345 ( .x(n3122), .a(n662), .b(n1380), .c(n1398) );
	aoi22_1 U2346 ( .x(n3029), .a(n1095), .b(n1380), .c(n1197), .d(n594) );
	and4i_5 U2347 ( .x(n840), .a(n841), .b(n2334), .c(n3758), .d(n3753) );
	inv_16 U2348 ( .x(___cell__39620_net143962), .a(Imm[16]) );
	inv_10 U2349 ( .x(n1334), .a(n3475) );
	nand2i_2 U235 ( .x(n3924), .a(n718), .b(n2783) );
	oai22_2 U2350 ( .x(n2116), .a(n884), .b(n1616), .c(___cell__39620_net143658),
		.d(n2112) );
	nor2i_3 U2351 ( .x(n1094), .a(n1095), .b(n884) );
	aoi22_1 U2352 ( .x(n2801), .a(n544), .b(___cell__39620_net143864), .c(n1204),
		.d(n2803) );
	aoi221_1 U2353 ( .x(n2580), .a(n2581), .b(n1267), .c(reg_out_B[25]), .d(n1064),
		.e(n2582) );
	aoi222_2 U2354 ( .x(n2182), .a(n1256), .b(n1999), .c(n2183), .d(n2184),
		.e(n2185), .f(n636) );
	inv_14 U2355 ( .x(n1256), .a(n1634) );
	nand2_5 U2356 ( .x(n1622), .a(n923), .b(net149167) );
	inv_1 U2357 ( .x(n632), .a(Imm[18]) );
	nor2_0 U2358 ( .x(n801), .a(IR_opcode_field[2]), .b(IR_opcode_field[4]) );
	nand2i_0 U2359 ( .x(n1614), .a(IR_opcode_field[4]), .b(IR_opcode_field[5]) );
	nand2i_2 U236 ( .x(n3925), .a(n4008), .b(n2784) );
	buf_10 U2360 ( .x(n634), .a(reg_out_A[23]) );
	inv_0 U2361 ( .x(n641), .a(Imm[6]) );
	inv_2 U2362 ( .x(n642), .a(n641) );
	exnor2_1 U2363 ( .x(n1502), .a(reg_out_B[17]), .b(n902) );
	aoi22_1 U2364 ( .x(n2928), .a(reg_out_B[17]), .b(n2929), .c(n2024), .d(n2930) );
	nand3i_4 U2365 ( .x(n646), .a(___cell__39620_net144175), .b(n1528), .c(n645) );
	inv_2 U2366 ( .x(n645), .a(n1524) );
	nor2_8 U2367 ( .x(n777), .a(Imm[20]), .b(n631) );
	nor2i_3 U2368 ( .x(n651), .a(n896), .b(n1573) );
	or3i_3 U2369 ( .x(n789), .a(N1729), .b(___cell__39620_net147731), .c(___cell__39620_net143660) );
	exnor2_1 U237 ( .x(n1503), .a(reg_out_B[16]), .b(n893) );
	inv_2 U2370 ( .x(n652), .a(___cell__39620_net144360) );
	nand4_1 U2371 ( .x(n1548), .a(n1954), .b(n653), .c(n1953), .d(n1952) );
	ao221_4 U2372 ( .x(n2939), .a(n3902), .b(n654), .c(n3903), .d(n655), .e(n516) );
	inv_0 U2373 ( .x(n654), .a(n621) );
	inv_2 U2374 ( .x(n655), .a(___cell__39620_net144406) );
	inv_2 U2375 ( .x(n656), .a(reg_out_B[31]) );
	nand2i_8 U2376 ( .x(n1700), .a(n766), .b(n1701) );
	nand2_8 U2377 ( .x(n1633), .a(n896), .b(reg_out_B[4]) );
	oai221_5 U2378 ( .x(n2600), .a(n1324), .b(n4005), .c(n3421), .d(n4006),
		.e(n1806) );
	inv_2 U2379 ( .x(n657), .a(n947) );
	inv_14 U238 ( .x(n631), .a(___cell__39620_net143962) );
	nand2i_6 U2380 ( .x(n1688), .a(reg_out_B[3]), .b(n1689) );
	and2_8 U2381 ( .x(n658), .a(n1689), .b(reg_out_A[30]) );
	oai211_2 U2382 ( .x(n4061), .a(___cell__39620_net143287), .b(n966), .c(n967),
		.d(n968) );
	inv_0 U2383 ( .x(n659), .a(reg_out_B[3]) );
	oai211_2 U2384 ( .x(n4056), .a(___cell__39620_net143287), .b(n957), .c(n958),
		.d(n959) );
	inv_6 U2385 ( .x(n660), .a(n3071) );
	nand2i_8 U2386 ( .x(n1642), .a(reg_out_B[2]), .b(n882) );
	oai211_2 U2387 ( .x(n1968), .a(n855), .b(n3596), .c(n1040), .d(n3353) );
	inv_16 U2388 ( .x(n815), .a(n828) );
	ao31_4 U2389 ( .x(n2402), .a(n2629), .b(n763), .c(n828), .d(n819) );
	inv_2 U239 ( .x(n1861), .a(N1748) );
	ao22_1 U2390 ( .x(n3378), .a(n828), .b(n3307), .c(n826), .d(n813) );
	nand2_2 U2391 ( .x(n1419), .a(n664), .b(___cell__39620_net144328) );
	nand2_8 U2392 ( .x(n665), .a(n664), .b(___cell__39620_net144328) );
	inv_16 U2393 ( .x(___cell__39620_net144328), .a(___cell__39620_net144324) );
	inv_2 U2394 ( .x(___cell__39620_net144326), .a(net151578) );
	oai221_2 U2395 ( .x(n2874), .a(n752), .b(n1635), .c(n3447), .d(n4009),
		.e(n2850) );
	inv_14 U2396 ( .x(n1728), .a(n1159) );
	oai22_2 U2397 ( .x(n3382), .a(n1580), .b(n915), .c(n1578), .d(n1642) );
	oa22_2 U2398 ( .x(n761), .a(n1570), .b(n1631), .c(___cell__39620_net144257),
		.d(n4012) );
	inv_3 U2399 ( .x(n833), .a(reg_out_A[4]) );
	nand2i_5 U240 ( .x(n3764), .a(n751), .b(n3763) );
	nor2i_3 U2400 ( .x(n666), .a(n667), .b(___cell__39620_net144329) );
	inv_4 U2401 ( .x(n1624), .a(n666) );
	inv_0 U2402 ( .x(n667), .a(___cell__39620_net144331) );
	ao22_3 U2403 ( .x(n3166), .a(n3981), .b(n668), .c(n766), .d(n818) );
	inv_2 U2404 ( .x(n668), .a(n670) );
	nand2_2 U2405 ( .x(n1637), .a(n669), .b(n1638) );
	inv_1 U2406 ( .x(n669), .a(___cell__39620_net144175) );
	nand2_5 U2407 ( .x(n670), .a(n669), .b(n1638) );
	nand3_2 U2408 ( .x(n3007), .a(n3011), .b(n515), .c(n3015) );
	nand2i_8 U2409 ( .x(___cell__39620_net144329), .a(Imm[5]), .b(n773) );
	inv_4 U241 ( .x(n3639), .a(n3638) );
	nand2i_2 U2410 ( .x(n3948), .a(n1632), .b(n525) );
	nand3_4 U2411 ( .x(n2299), .a(N1861), .b(n4000), .c(___cell__39620_net147732) );
	aoi22_1 U2412 ( .x(n3191), .a(N1831), .b(n4000), .c(N1964), .d(___cell__39620_net145508) );
	or2_8 U2413 ( .x(n3628), .a(n3395), .b(n610) );
	inv_3 U2414 ( .x(n3395), .a(n3626) );
	nor2_0 U2415 ( .x(___cell__39620_net143982), .a(___cell__39620_net143693),
		.b(___cell__39620_net143983) );
	nor2_3 U2418 ( .x(n1962), .a(reg_out_B[16]), .b(reg_out_B[17]) );
	inv_0 U2419 ( .x(n1866), .a(reg_out_B[16]) );
	nand2i_4 U242 ( .x(n2722), .a(n751), .b(n3818) );
	or2_8 U2420 ( .x(n3511), .a(n1072), .b(n672) );
	and2_8 U2421 ( .x(n673), .a(net149167), .b(n891) );
	nand2i_2 U2422 ( .x(n1072), .a(net149167), .b(n891) );
	inv_16 U2423 ( .x(n1289), .a(n1607) );
	oai21_6 U2424 ( .x(n2384), .a(n3524), .b(n4005), .c(n3572) );
	nand2i_2 U2425 ( .x(n3572), .a(n4140), .b(n1043) );
	and3i_4 U2426 ( .x(n674), .a(___cell__39620_net147731), .b(n676), .c(n514) );
	inv_12 U2427 ( .x(n784), .a(n674) );
	and2_8 U2428 ( .x(n676), .a(n677), .b(___cell__39620_net144344) );
	inv_0 U2429 ( .x(n677), .a(IR_opcode_field[0]) );
	nand2i_2 U243 ( .x(n3884), .a(n4005), .b(n3658) );
	or2_8 U2430 ( .x(n3646), .a(n3497), .b(n610) );
	inv_3 U2431 ( .x(n3497), .a(n3645) );
	inv_16 U2432 ( .x(n942), .a(n941) );
	mux2i_3 U2433 ( .x(n2710), .d0(n3536), .sl(net149120), .d1(n510) );
	inv_10 U2434 ( .x(n3536), .a(n3535) );
	nor2i_3 U2435 ( .x(n1663), .a(n2006), .b(n1543) );
	oai22_3 U2436 ( .x(n2570), .a(n1573), .b(n890), .c(___cell__39620_net144257),
		.d(n1651) );
	inv_16 U2437 ( .x(n1651), .a(n811) );
	inv_0 U2438 ( .x(___cell__39620_net144605), .a(Imm[29]) );
	buf_16 U2439 ( .x(n832), .a(reg_out_A[1]) );
	nand2i_6 U244 ( .x(n3658), .a(n3542), .b(n3627) );
	buf_16 U2440 ( .x(n921), .a(n937) );
	inv_14 U2441 ( .x(n681), .a(n680) );
	aoi22_2 U2442 ( .x(n3114), .a(n502), .b(n3116), .c(n3117), .d(___cell__39620_net143722) );
	mux2i_2 U2443 ( .x(n3117), .d0(n3417), .sl(n816), .d1(n3358) );
	nand2i_2 U2444 ( .x(n2975), .a(n621), .b(n3010) );
	aoi22_2 U2445 ( .x(n1967), .a(n1964), .b(n1968), .c(n1330), .d(n1969) );
	aoi22_2 U2446 ( .x(n3021), .a(n1971), .b(n3022), .c(n1330), .d(n1968) );
	nand4_1 U2447 ( .x(n3010), .a(n3921), .b(n3920), .c(n3919), .d(n3918) );
	exnor2_1 U2448 ( .x(n1476), .a(reg_out_A[29]), .b(reg_out_B[29]) );
	inv_10 U2449 ( .x(n747), .a(n685) );
	inv_5 U245 ( .x(n3306), .a(n3303) );
	nand2i_8 U2450 ( .x(n1557), .a(n1039), .b(n1558) );
	buf_12 U2451 ( .x(n686), .a(reg_out_A[22]) );
	nor2i_3 U2452 ( .x(n1134), .a(n838), .b(n1122) );
	nor2i_3 U2453 ( .x(n1133), .a(n838), .b(n1120) );
	aoai211_1 U2454 ( .x(n2790), .a(n749), .b(n530), .c(n1064), .d(reg_out_B[20]) );
	exnor2_1 U2455 ( .x(n1493), .a(reg_out_B[20]), .b(n749) );
	inv_16 U2456 ( .x(n691), .a(n940) );
	inv_16 U2457 ( .x(n692), .a(n691) );
	nand2_6 U2458 ( .x(n3303), .a(n3304), .b(n3305) );
	nand2_2 U2459 ( .x(n3647), .a(n923), .b(n634) );
	nand2i_2 U246 ( .x(n3885), .a(n1625), .b(n3303) );
	or3i_2 U2461 ( .x(n1940), .a(n2002), .b(n693), .c(n1521) );
	inv_0 U2462 ( .x(n693), .a(IR_function_field[4]) );
	ao22_6 U2463 ( .x(n1996), .a(reg_out_A[20]), .b(n3575), .c(n3464), .d(n799) );
	buf_16 U2464 ( .x(n694), .a(net149107) );
	nand2_8 U2465 ( .x(n696), .a(n713), .b(n928) );
	ao211_5 U2466 ( .x(n2857), .a(n3374), .b(n625), .c(n698), .d(n697) );
	and2_2 U2467 ( .x(n698), .a(n699), .b(n2995) );
	inv_2 U2468 ( .x(n699), .a(n727) );
	inv_16 U2469 ( .x(n816), .a(n879) );
	nand2i_2 U247 ( .x(n3886), .a(___cell__39620_net144062), .b(n3034) );
	inv_0 U2470 ( .x(n700), .a(n702) );
	nand2_8 U2471 ( .x(n703), .a(n701), .b(n1661) );
	nand2i_5 U2472 ( .x(n3613), .a(n3612), .b(n3598) );
	nand2i_2 U2473 ( .x(n3499), .a(n1647), .b(n1689) );
	oa22_2 U2474 ( .x(n856), .a(n815), .b(n761), .c(n1573), .d(n915) );
	inv_16 U2475 ( .x(n901), .a(n900) );
	or3i_4 U2476 ( .x(n704), .a(N1663), .b(n705), .c(___cell__39620_net143872) );
	inv_0 U2477 ( .x(n705), .a(___cell__39620_net147732) );
	inv_16 U2478 ( .x(n809), .a(n706) );
	inv_2 U2479 ( .x(n707), .a(n808) );
	nand2i_2 U248 ( .x(n3904), .a(n1562), .b(n2719) );
	inv_0 U2480 ( .x(n710), .a(IR_opcode_field[3]) );
	aoi21_1 U2481 ( .x(n802), .a(IR_opcode_field[0]), .b(___cell__39620_net143655),
		.c(n800) );
	nand2i_0 U2482 ( .x(n808), .a(IR_opcode_field[1]), .b(n810) );
	inv_2 U2483 ( .x(n726), .a(n816) );
	inv_5 U2484 ( .x(n1451), .a(n816) );
	nand2i_6 U2485 ( .x(n3619), .a(n3618), .b(n3598) );
	inv_2 U2486 ( .x(n841), .a(n3759) );
	nand2i_2 U2487 ( .x(n3906), .a(n4004), .b(n3610) );
	nand4_1 U2488 ( .x(n1000), .a(n3699), .b(n2153), .c(n2146), .d(n2158) );
	nand2i_2 U2489 ( .x(n2158), .a(n1692), .b(n2837) );
	inv_5 U249 ( .x(n1971), .a(n1562) );
	and4i_2 U2490 ( .x(n2153), .a(n2149), .b(n2154), .c(n2155), .d(n2156) );
	oai22_6 U2491 ( .x(n3384), .a(n1564), .b(n915), .c(n1219), .d(n1642) );
	inv_10 U2492 ( .x(n902), .a(n862) );
	ao21_4 U2493 ( .x(n3963), .a(n3415), .b(n711), .c(n712) );
	inv_0 U2494 ( .x(n711), .a(n1451) );
	inv_16 U2495 ( .x(n908), .a(n907) );
	inv_16 U2496 ( .x(n907), .a(reg_out_A[10]) );
	inv_16 U2497 ( .x(n3598), .a(n1557) );
	inv_4 U2498 ( .x(n714), .a(n1067) );
	inv_2 U2499 ( .x(n715), .a(___cell__39620_net144374) );
	buf_1 U25 ( .x(n635), .a(reg_out_A[23]) );
	nand2i_2 U250 ( .x(n3905), .a(n1565), .b(n3613) );
	nand2i_8 U2500 ( .x(___cell__39620_net144062), .a(n891), .b(n717) );
	or2_4 U2501 ( .x(___cell__39620_net144374), .a(n637), .b(n717) );
	or2_4 U2502 ( .x(n719), .a(n637), .b(n717) );
	or2_4 U2503 ( .x(n718), .a(n637), .b(n717) );
	inv_5 U2504 ( .x(n3452), .a(n3451) );
	aoi221_5 U2505 ( .x(n720), .a(n2133), .b(n723), .c(n722), .d(n721), .e(n724) );
	inv_2 U2506 ( .x(n721), .a(n727) );
	inv_2 U2507 ( .x(n723), .a(n1635) );
	ao22_3 U2508 ( .x(n724), .a(n1249), .b(n1997), .c(n1256), .d(n847) );
	nand2_1 U2509 ( .x(n727), .a(n726), .b(n725) );
	nand2i_4 U251 ( .x(n3059), .a(n3585), .b(n3817) );
	nor2i_3 U2510 ( .x(n728), .a(n725), .b(n726) );
	inv_10 U2511 ( .x(n1635), .a(n728) );
	inv_5 U2512 ( .x(n3317), .a(n2233) );
	oai22_4 U2513 ( .x(n2130), .a(n3504), .b(n536), .c(n1577), .d(n1629) );
	inv_2 U2514 ( .x(n1178), .a(n3327) );
	inv_16 U2515 ( .x(n887), .a(n886) );
	nand2_1 U2516 ( .x(n3327), .a(n3328), .b(n3329) );
	oai21_5 U2517 ( .x(n3410), .a(n3411), .b(n815), .c(n3412) );
	oai211_2 U2518 ( .x(n4059), .a(n963), .b(___cell__39620_net147731), .c(n964),
		.d(n965) );
	and4i_2 U2519 ( .x(n963), .a(n1413), .b(n1410), .c(n1411), .d(n1412) );
	nand2i_2 U252 ( .x(n3301), .a(n1563), .b(n926) );
	inv_2 U2520 ( .x(n729), .a(n816) );
	oai221_2 U2522 ( .x(n3903), .a(n752), .b(n1636), .c(n3411), .d(n1632),
		.e(n2925) );
	aoi22_2 U2523 ( .x(n2891), .a(n910), .b(n2892), .c(n2024), .d(n2857) );
	and2_8 U2524 ( .x(n735), .a(___cell__39620_net144356), .b(___cell__39620_net143655) );
	inv_14 U2525 ( .x(n946), .a(n735) );
	inv_4 U2526 ( .x(___cell__39620_net143655), .a(n804) );
	nor2_1 U2527 ( .x(___cell__39620_net144356), .a(n805), .b(___cell__39620_net144166) );
	oai22_6 U2528 ( .x(n2888), .a(n1586), .b(n881), .c(n822), .d(n1654) );
	inv_10 U2529 ( .x(n773), .a(n771) );
	inv_5 U2530 ( .x(n1257), .a(n2690) );
	oai211_2 U2531 ( .x(n3289), .a(n3434), .b(n1560), .c(n1040), .d(n2810) );
	ao22_6 U2532 ( .x(n2133), .a(n3336), .b(n812), .c(reg_out_A[20]), .d(n3584) );
	inv_3 U2533 ( .x(n3334), .a(n3336) );
	nand2_2 U2534 ( .x(n3336), .a(n3337), .b(n3338) );
	nor2_8 U2535 ( .x(n813), .a(n1560), .b(n825) );
	oai22_3 U2536 ( .x(n3545), .a(n915), .b(n1646), .c(n1642), .d(n1644) );
	oai22_3 U2537 ( .x(n2236), .a(n1642), .b(n1649), .c(n915), .d(n1647) );
	nor2i_8 U2538 ( .x(n737), .a(n768), .b(n825) );
	inv_16 U2539 ( .x(n883), .a(n825) );
	nand2i_2 U254 ( .x(n3296), .a(n1654), .b(n874) );
	or2_4 U2540 ( .x(n4009), .a(n816), .b(n815) );
	nand2i_8 U2541 ( .x(n1558), .a(n855), .b(n1728) );
	inv_10 U2542 ( .x(n1283), .a(n3467) );
	inv_0 U2543 ( .x(n739), .a(n816) );
	inv_12 U2544 ( .x(n3313), .a(n3312) );
	oai22_5 U2545 ( .x(n2995), .a(n1587), .b(n822), .c(n1583), .d(n881) );
	aoi22_1 U2546 ( .x(n2431), .a(n2432), .b(n590), .c(n1249), .d(n2433) );
	nand2i_2 U2547 ( .x(n3930), .a(n4009), .b(n2690) );
	aoi22_2 U2548 ( .x(n2044), .a(n1683), .b(n2045), .c(___cell__39620_net144517),
		.d(n1995) );
	oai22_4 U2549 ( .x(n2045), .a(n1577), .b(n871), .c(n500), .d(n4125) );
	nand2i_2 U255 ( .x(n3892), .a(n4008), .b(n2991) );
	aoai211_5 U2550 ( .x(n740), .a(n3862), .b(n741), .c(n742), .d(n1444) );
	inv_5 U2551 ( .x(n1449), .a(n740) );
	inv_2 U2552 ( .x(n741), .a(n1451) );
	nand4i_2 U2553 ( .x(n3862), .a(n1278), .b(n3860), .c(n2807), .d(n3412) );
	nand2i_1 U2554 ( .x(n3759), .a(n1608), .b(n3321) );
	nand2_0 U2555 ( .x(n2912), .a(n640), .b(n902) );
	exnor2_1 U2556 ( .x(n1501), .a(n902), .b(n640) );
	inv_0 U2557 ( .x(___cell__39620_net143954), .a(n640) );
	inv_16 U2558 ( .x(n745), .a(n744) );
	nand2i_2 U2559 ( .x(n2341), .a(n1632), .b(n1999) );
	nand2i_2 U256 ( .x(n3894), .a(n4010), .b(n2992) );
	aoi22_1 U2560 ( .x(n1998), .a(n1999), .b(n504), .c(n1256), .d(n2000) );
	mux2_4 U2561 ( .x(n746), .d0(n3546), .sl(n816), .d1(n3442) );
	aoi221_1 U2562 ( .x(n2188), .a(n2189), .b(___cell__39620_net144345), .c(n912),
		.d(n2190), .e(n1130) );
	inv_2 U2563 ( .x(n3604), .a(n3491) );
	nor2i_0 U2564 ( .x(n2161), .a(net151578), .b(n1656) );
	exnor2_1 U2565 ( .x(n1465), .a(n912), .b(net151578) );
	inv_16 U2566 ( .x(n749), .a(n748) );
	nor2_3 U2567 ( .x(n2146), .a(n2143), .b(n2141) );
	buf_5 U2568 ( .x(n750), .a(n2236) );
	and4i_3 U2569 ( .x(n1262), .a(n2773), .b(n2775), .c(n2776), .d(n2777) );
	exnor2_1 U257 ( .x(n1491), .a(n628), .b(n566) );
	or2_8 U2570 ( .x(n1281), .a(n1684), .b(n671) );
	nand2i_3 U2571 ( .x(n1684), .a(net149167), .b(n1685) );
	inv_4 U2572 ( .x(n1772), .a(N333) );
	oai22_2 U2574 ( .x(n2773), .a(n2774), .b(n1616), .c(n865), .d(n1166) );
	oa211_5 U2575 ( .x(n865), .a(n3629), .b(n1043), .c(n2765), .d(n3859) );
	nand2i_1 U2576 ( .x(n3603), .a(n1587), .b(n896) );
	nand2i_1 U2577 ( .x(n3607), .a(n1219), .b(n896) );
	nand2i_2 U2578 ( .x(n3608), .a(n1564), .b(n896) );
	nand2i_2 U2579 ( .x(n1672), .a(n1673), .b(n896) );
	nand2i_2 U258 ( .x(n3528), .a(n891), .b(n2992) );
	nand2i_3 U2580 ( .x(n3596), .a(___cell__39620_net144257), .b(n896) );
	oa21_6 U2581 ( .x(n752), .a(n2475), .b(reg_out_B[3]), .c(n3551) );
	nand2i_4 U2582 ( .x(n3551), .a(n1648), .b(n3584) );
	inv_16 U2583 ( .x(n753), .a(___cell__39620_net144655) );
	and2_8 U2584 ( .x(n754), .a(n839), .b(reg_out_B[3]) );
	inv_16 U2585 ( .x(n1629), .a(n754) );
	aoi22_1 U2586 ( .x(n2479), .a(n2435), .b(n2277), .c(n2436), .d(n914) );
	aoi21_1 U2587 ( .x(n1082), .a(n914), .b(n530), .c(n1064) );
	aoi22_1 U2588 ( .x(n2281), .a(n2268), .b(n894), .c(n823), .d(n914) );
	inv_2 U2589 ( .x(n1648), .a(n914) );
	nand2i_5 U259 ( .x(n3375), .a(n1219), .b(n3592) );
	aoi22_1 U2590 ( .x(n2562), .a(n2266), .b(n914), .c(n1391), .d(n4134) );
	exnor2_1 U2591 ( .x(n1459), .a(reg_out_B[8]), .b(n914) );
	inv_16 U2592 ( .x(n2475), .a(n2283) );
	inv_0 U2593 ( .x(n755), .a(n703) );
	inv_2 U2594 ( .x(n756), .a(n1658) );
	inv_12 U2595 ( .x(n1249), .a(n1632) );
	inv_0 U2596 ( .x(n757), .a(n784) );
	inv_0 U2597 ( .x(n758), .a(___cell__39620_net144406) );
	and3i_1 U2598 ( .x(n760), .a(reg_out_B[4]), .b(n759), .c(n1552) );
	inv_0 U2599 ( .x(n899), .a(n760) );
	inv_8 U26 ( .x(n1654), .a(reg_out_A[3]) );
	inv_8 U260 ( .x(n529), .a(n1629) );
	inv_3 U2600 ( .x(n1570), .a(n583) );
	oai211_3 U2601 ( .x(n2789), .a(n2655), .b(n1186), .c(n2785), .d(n2790) );
	ao21_4 U2602 ( .x(n3415), .a(n2888), .b(n828), .c(n762) );
	inv_0 U2604 ( .x(n763), .a(reg_out_B[3]) );
	inv_0 U2605 ( .x(n764), .a(n621) );
	inv_2 U2606 ( .x(n765), .a(n670) );
	nand2i_4 U2607 ( .x(n2296), .a(n1592), .b(N338) );
	inv_16 U2608 ( .x(N3304), .a(___cell__6067_net21981) );
	and3i_4 U2609 ( .x(n964), .a(n3165), .b(n3983), .c(n3164) );
	inv_5 U261 ( .x(n1250), .a(n2851) );
	ao222_4 U2610 ( .x(n2930), .a(reg_out_B[1]), .b(n3365), .c(n827), .d(n767),
		.e(n3036), .f(n768) );
	inv_2 U2611 ( .x(n767), .a(n1634) );
	inv_2 U2612 ( .x(n768), .a(n4009) );
	nor3_3 U2613 ( .x(n982), .a(n2662), .b(n2669), .c(n2666) );
	inv_2 U2614 ( .x(net150643), .a(___cell__39620_net143767) );
	nor2_0 U2615 ( .x(___cell__39620_net143767), .a(n4140), .b(n770) );
	inv_16 U2616 ( .x(___cell__39620_net147732), .a(___cell__39620_net147731) );
	nand2i_6 U2618 ( .x(___cell__39620_net144324), .a(N69), .b(n773) );
	nor2_1 U2619 ( .x(___cell__39620_net145077), .a(Imm[14]), .b(Imm[11]) );
	nand2i_2 U262 ( .x(n3373), .a(n1644), .b(n874) );
	nand2i_4 U2620 ( .x(n778), .a(Imm[17]), .b(n777) );
	oai221_4 U2621 ( .x(n790), .a(n792), .b(___cell__39620_net144406), .c(n793),
		.d(n784), .e(n791) );
	inv_6 U2622 ( .x(n793), .a(___cell__39620_net147278) );
	oai211_3 U2623 ( .x(n788), .a(n503), .b(n785), .c(n787), .d(n789) );
	aoi23_4 U2624 ( .x(n787), .a(n786), .b(___cell__39620_net147732), .c(N1762),
		.d(___cell__39620_net143326), .e(___cell__39620_net145150) );
	nor2i_5 U2625 ( .x(n786), .a(net151622), .b(n734) );
	inv_16 U2626 ( .x(___cell__39620_net145150), .a(___cell__39620_net143710) );
	nand2i_4 U2627 ( .x(n785), .a(___cell__39620_net144343), .b(___cell__39620_net143326) );
	nor2i_5 U2628 ( .x(___cell__39620_net143784), .a(___cell__39620_net143785),
		.b(n503) );
	nand4i_4 U2629 ( .x(___cell__39620_net145427), .a(___cell__39620_net145428),
		.b(___cell__39620_net145429), .c(n796), .d(n797) );
	nand2i_2 U263 ( .x(n3377), .a(n1655), .b(n874) );
	inv_16 U2630 ( .x(___cell__39620_net145508), .a(___cell__39620_net143845) );
	nand3i_5 U2631 ( .x(n796), .a(___cell__39620_net144062), .b(___cell__39620_net147296),
		.c(n798) );
	nand2i_6 U2632 ( .x(n794), .a(n4140), .b(n795) );
	inv_16 U2633 ( .x(net151904), .a(___cell__39620_net144331) );
	inv_16 U2634 ( .x(___cell__39620_net144331), .a(Imm[4]) );
	inv_10 U2635 ( .x(n803), .a(IR_opcode_field[2]) );
	and2_5 U2636 ( .x(___cell__39620_net145037), .a(n803), .b(net151497) );
	nand2i_8 U2637 ( .x(___cell__39620_net143710), .a(n803), .b(___cell__39620_net144309) );
	and3i_1 U2638 ( .x(n800), .a(___cell__39620_net143653), .b(n801), .c(IR_opcode_field[5]) );
	or3i_1 U2639 ( .x(n804), .a(IR_opcode_field[5]), .b(IR_opcode_field[4]),
		.c(IR_opcode_field[1]) );
	oai22_5 U264 ( .x(n2690), .a(n1585), .b(n881), .c(n1629), .d(n1655) );
	nand2i_8 U2640 ( .x(___cell__39620_net147731), .a(n807), .b(N3304) );
	nand2i_8 U2641 ( .x(___cell__39620_net143287), .a(n568), .b(N3304) );
	nand2i_6 U2642 ( .x(___cell__39620_net144199), .a(___cell__39620_net144200),
		.b(n708) );
	nand2_8 U2643 ( .x(___cell__39620_net143658), .a(___cell__39620_net144303),
		.b(n708) );
	buf_2 U2644 ( .x(n926), .a(n531) );
	inv_16 U2645 ( .x(n1602), .a(Imm[2]) );
	inv_2 U2646 ( .x(net149616), .a(Imm[9]) );
	nand2i_0 U2647 ( .x(n1535), .a(IR_function_field[0]), .b(IR_function_field[1]) );
	inv_2 U2648 ( .x(n1534), .a(IR_function_field[1]) );
	ao22_6 U2649 ( .x(n2000), .a(n3346), .b(n812), .c(n628), .d(n3584) );
	nand2i_3 U265 ( .x(n3394), .a(n3395), .b(n3396) );
	inv_0 U2650 ( .x(n812), .a(reg_out_B[3]) );
	inv_4 U2651 ( .x(n3345), .a(n3346) );
	nand2_2 U2652 ( .x(n3346), .a(n3347), .b(n3348) );
	inv_3 U2653 ( .x(n1560), .a(n815) );
	inv_2 U2654 ( .x(n814), .a(n1569) );
	nand2_2 U2655 ( .x(n3318), .a(n3319), .b(n3320) );
	mux2_4 U2656 ( .x(n870), .d0(n3446), .sl(n694), .d1(n589) );
	and2_3 U2657 ( .x(n1978), .a(n817), .b(n905) );
	aoi211_1 U2658 ( .x(n2127), .a(n2079), .b(n2128), .c(n1108), .d(n1109) );
	inv_5 U266 ( .x(n3391), .a(n3496) );
	inv_2 U2660 ( .x(n818), .a(n817) );
	nand2i_0 U2661 ( .x(n2297), .a(n4039), .b(n3057) );
	oai21_3 U2662 ( .x(n3760), .a(net149122), .b(n840), .c(n2336) );
	inv_0 U2663 ( .x(n819), .a(n1159) );
	inv_2 U2664 ( .x(n820), .a(n819) );
	nand2i_2 U2665 ( .x(n3881), .a(n4003), .b(n3599) );
	oai22_1 U2666 ( .x(n2330), .a(n1087), .b(n4038), .c(___cell__39620_net143693),
		.d(___cell__39620_net144572) );
	and4_5 U2667 ( .x(n2314), .a(n2313), .b(n2316), .c(n2315), .d(n821) );
	nand2i_0 U2668 ( .x(n2315), .a(n4140), .b(n1318) );
	nand2i_3 U2669 ( .x(n3599), .a(n3597), .b(n3598) );
	buf_16 U2670 ( .x(n822), .a(n4012) );
	nor2_3 U2671 ( .x(n823), .a(n1688), .b(n824) );
	inv_0 U2672 ( .x(n824), .a(n815) );
	nand3_5 U2673 ( .x(n3702), .a(n2186), .b(n3701), .c(n2182) );
	buf_16 U2675 ( .x(net149120), .a(net149107) );
	oai21_1 U2677 ( .x(n3247), .a(n3237), .b(n3238), .c(n943) );
	oai21_1 U2678 ( .x(n3241), .a(n943), .b(___cell__39620_net144199), .c(n1618) );
	nor3_0 U2679 ( .x(n3256), .a(n1521), .b(IR_function_field[2]), .c(IR_function_field[4]) );
	inv_2 U2680 ( .x(n826), .a(n1573) );
	inv_10 U2681 ( .x(n829), .a(n830) );
	inv_6 U2682 ( .x(n909), .a(reg_out_A[18]) );
	exnor2_1 U2684 ( .x(n1513), .a(reg_out_B[11]), .b(n901) );
	inv_0 U2685 ( .x(n1907), .a(reg_out_B[11]) );
	inv_10 U2686 ( .x(net149628), .a(net149627) );
	nand2i_1 U2687 ( .x(n3640), .a(n1603), .b(n902) );
	aoi21_1 U2688 ( .x(n2369), .a(n885), .b(n1733), .c(n1179) );
	aoi21_1 U2689 ( .x(n2147), .a(n885), .b(n2148), .c(n1117) );
	inv_16 U269 ( .x(n874), .a(n1622) );
	aoai211_1 U2690 ( .x(n2357), .a(n885), .b(n530), .c(n1064), .d(n536) );
	exnor2_1 U2691 ( .x(n1473), .a(net149167), .b(n885) );
	exnor2_1 U2692 ( .x(n1474), .a(reg_out_B[3]), .b(n885) );
	inv_0 U2693 ( .x(___cell__39620_net143720), .a(Imm[7]) );
	inv_0 U2694 ( .x(___cell__39620_net144572), .a(Imm[30]) );
	aoi22_2 U2695 ( .x(n2709), .a(n2710), .b(n1267), .c(n2711), .d(n502) );
	inv_2 U2696 ( .x(net151577), .a(Imm[5]) );
	mux2i_1 U2697 ( .x(n1951), .d0(n1446), .sl(reg_out_B[0]), .d1(n1527) );
	exnor2_1 U2698 ( .x(n3274), .a(reg_out_B[0]), .b(n942) );
	nand2i_0 U2699 ( .x(n1628), .a(IR_function_field[0]), .b(reg_out_B[0]) );
	inv_8 U27 ( .x(___cell__39620_net143983), .a(Imm[15]) );
	nand2i_2 U270 ( .x(n3461), .a(n1563), .b(n874) );
	nand2_0 U2700 ( .x(n1568), .a(reg_out_B[0]), .b(IR_function_field[0]) );
	nor2i_0 U2701 ( .x(n2001), .a(reg_out_B[0]), .b(n1524) );
	nand2i_0 U2702 ( .x(n1659), .a(reg_out_B[0]), .b(n645) );
	nand2_0 U2703 ( .x(n3257), .a(IR_function_field[3]), .b(IR_function_field[1]) );
	or3i_2 U2704 ( .x(n1538), .a(IR_function_field[2]), .b(IR_function_field[4]),
		.c(IR_function_field[3]) );
	nand2_0 U2705 ( .x(n2588), .a(Imm[24]), .b(n541) );
	exnor2_1 U2706 ( .x(n1486), .a(n541), .b(Imm[24]) );
	aoi21_1 U2707 ( .x(n1104), .a(n852), .b(n530), .c(n1064) );
	nor2i_3 U2708 ( .x(n1092), .a(n852), .b(n1093) );
	nor2i_3 U2709 ( .x(n1119), .a(n852), .b(n1120) );
	nand2i_2 U271 ( .x(n3494), .a(n1654), .b(n1689) );
	nor2i_3 U2710 ( .x(n1088), .a(n852), .b(n695) );
	nor2i_3 U2711 ( .x(n1121), .a(n852), .b(n1122) );
	exnor2_1 U2712 ( .x(n1461), .a(n4146), .b(n852) );
	inv_2 U2713 ( .x(n1655), .a(reg_out_A[7]) );
	exnor2_1 U2714 ( .x(n1462), .a(Imm[7]), .b(n852) );
	nand2_0 U2715 ( .x(n2068), .a(n852), .b(Imm[7]) );
	ao21_6 U2716 ( .x(n3741), .a(n861), .b(n835), .c(n1728) );
	nand2i_2 U2717 ( .x(n3645), .a(n925), .b(n887) );
	nand2i_2 U2718 ( .x(n3637), .a(n925), .b(n628) );
	nand2i_2 U2719 ( .x(n3654), .a(n925), .b(n686) );
	and2_3 U272 ( .x(n506), .a(n3494), .b(n3495) );
	nand2i_2 U2720 ( .x(n3588), .a(n925), .b(n894) );
	nand2i_2 U2721 ( .x(n3626), .a(n925), .b(n749) );
	nand2i_2 U2722 ( .x(n3664), .a(n925), .b(n914) );
	nand2i_4 U2723 ( .x(n3577), .a(n925), .b(n609) );
	nand2i_2 U2724 ( .x(n3589), .a(n925), .b(n908) );
	oai21_2 U2725 ( .x(n1834), .a(n1646), .b(n890), .c(n1835) );
	aoi22_1 U2726 ( .x(n2907), .a(reg_out_B[18]), .b(n1064), .c(n633), .d(___cell__39620_net145617) );
	inv_0 U2727 ( .x(n1851), .a(reg_out_B[18]) );
	exnor2_1 U2728 ( .x(n1500), .a(n910), .b(reg_out_B[18]) );
	aoi22_1 U2729 ( .x(n2805), .a(___cell__39620_net144517), .b(n2806), .c(n1391),
		.d(n2045) );
	and2_3 U273 ( .x(n509), .a(n3490), .b(n3491) );
	aoi21_1 U2731 ( .x(n3213), .a(n3219), .b(n1267), .c(n3215) );
	inv_0 U2732 ( .x(n1532), .a(n4147) );
	exnor2_1 U2733 ( .x(n1457), .a(n4147), .b(n904) );
	aoi22_1 U2734 ( .x(n2873), .a(___cell__39620_net143722), .b(n2874), .c(___cell__39620_net143864),
		.d(n4129) );
	inv_0 U2736 ( .x(___cell__39620_net143694), .a(net149628) );
	nor2i_0 U2737 ( .x(n1227), .a(net149628), .b(___cell__39620_net143836) );
	exnor2_1 U2738 ( .x(n1460), .a(net149628), .b(n914) );
	nand2i_2 U2739 ( .x(n3488), .a(n1219), .b(n1685) );
	nand2_2 U274 ( .x(n2271), .a(n3308), .b(n3309) );
	nand2i_2 U2740 ( .x(n3566), .a(n1657), .b(n1685) );
	nand2i_2 U2741 ( .x(n3501), .a(n1647), .b(n1685) );
	nand2i_2 U2742 ( .x(n3487), .a(n1644), .b(n1685) );
	nand2i_2 U2743 ( .x(n3463), .a(___cell__39620_net144257), .b(n1685) );
	nand2i_1 U2744 ( .x(n3323), .a(n1587), .b(n1685) );
	nand2i_1 U2745 ( .x(n3472), .a(n1564), .b(n1685) );
	nand2i_1 U2746 ( .x(n3466), .a(n1580), .b(n1685) );
	nand2i_1 U2747 ( .x(n3543), .a(n1646), .b(n1685) );
	nand2i_2 U2748 ( .x(n3493), .a(n1655), .b(n1685) );
	nand2i_1 U2749 ( .x(n3469), .a(n1573), .b(n1685) );
	nand2i_2 U275 ( .x(n3387), .a(n1563), .b(n3584) );
	nand2i_1 U2750 ( .x(n3498), .a(n1654), .b(n1685) );
	nand2i_2 U2751 ( .x(n3396), .a(n1649), .b(n1685) );
	nand2i_2 U2752 ( .x(n3390), .a(n1656), .b(n1685) );
	nand2i_2 U2753 ( .x(n2729), .a(n1166), .b(n3856) );
	nand2i_4 U2754 ( .x(n995), .a(___cell__39620_net143287), .b(n3746) );
	inv_0 U2755 ( .x(net150830), .a(net149167) );
	inv_2 U2756 ( .x(n2177), .a(n2080) );
	nand2i_2 U2757 ( .x(n2355), .a(n1641), .b(n3760) );
	nand2_0 U2758 ( .x(n2018), .a(___cell__39620_net145617), .b(n4136) );
	nor2i_0 U2759 ( .x(n1212), .a(n4136), .b(___cell__39620_net143836) );
	inv_6 U276 ( .x(n3485), .a(n3483) );
	nor2i_0 U2760 ( .x(n1051), .a(n4136), .b(n1529) );
	exnor2_1 U2761 ( .x(n1458), .a(n904), .b(n4136) );
	inv_2 U2762 ( .x(n924), .a(n923) );
	oai22_2 U2763 ( .x(n2235), .a(n1649), .b(n889), .c(n1647), .d(n1651) );
	nand3i_0 U2764 ( .x(___cell__39620_net145419), .a(n2258), .b(___cell__39620_net147791),
		.c(___cell__39620_net143326) );
	inv_0 U2765 ( .x(net150620), .a(net149120) );
	inv_16 U2766 ( .x(n893), .a(n892) );
	oai211_2 U2767 ( .x(n4057), .a(n996), .b(___cell__39620_net147731), .c(n998),
		.d(n997) );
	nand2_1 U2768 ( .x(n3578), .a(n923), .b(n524) );
	inv_5 U2769 ( .x(n843), .a(n1971) );
	oai21_5 U277 ( .x(n3483), .a(net151904), .b(n1806), .c(n3484) );
	inv_4 U2770 ( .x(n2754), .a(n2711) );
	nor2i_8 U2771 ( .x(n844), .a(n3647), .b(n610) );
	nand2i_8 U2772 ( .x(n1604), .a(n1605), .b(n1606) );
	inv_0 U2773 ( .x(net150405), .a(net149122) );
	inv_4 U2774 ( .x(n846), .a(n2570) );
	oai22_2 U2775 ( .x(n847), .a(n1570), .b(n1629), .c(n512), .d(n536) );
	inv_16 U2776 ( .x(n3627), .a(n1604) );
	nand2i_2 U2777 ( .x(n3667), .a(n1632), .b(n847) );
	inv_0 U2778 ( .x(n848), .a(n816) );
	nor2_0 U2779 ( .x(n1158), .a(n820), .b(n1160) );
	aoi22_2 U278 ( .x(n853), .a(n858), .b(n883), .c(n855), .d(n854) );
	nor2_1 U2780 ( .x(n1185), .a(n820), .b(n1186) );
	inv_5 U2781 ( .x(n1749), .a(N369) );
	nand2i_2 U2782 ( .x(n3554), .a(n1578), .b(n1689) );
	nand2i_2 U2783 ( .x(n3473), .a(n1644), .b(n1689) );
	nand2i_1 U2784 ( .x(n3347), .a(n1564), .b(n1689) );
	nand2i_1 U2785 ( .x(n3337), .a(n1580), .b(n1689) );
	nand2i_2 U2786 ( .x(n3563), .a(n1657), .b(n1689) );
	nand2i_1 U2787 ( .x(n3404), .a(n1649), .b(n1689) );
	nand2i_1 U2788 ( .x(n3540), .a(n1646), .b(n1689) );
	nand2i_1 U2789 ( .x(n3328), .a(n1587), .b(n1689) );
	inv_10 U279 ( .x(n2067), .a(n1040) );
	nand2i_1 U2790 ( .x(n3319), .a(n1573), .b(n1689) );
	nand2i_2 U2791 ( .x(n3308), .a(n1656), .b(n1689) );
	nand2i_1 U2792 ( .x(n3490), .a(n1655), .b(n1689) );
	nand2_2 U2793 ( .x(n2333), .a(N337), .b(n2837) );
	inv_0 U2794 ( .x(n857), .a(reg_out_B[3]) );
	inv_2 U2795 ( .x(n858), .a(n1584) );
	inv_4 U2796 ( .x(n2083), .a(n2184) );
	inv_2 U2797 ( .x(n3383), .a(n3382) );
	and3i_3 U2798 ( .x(n994), .a(n2325), .b(n2333), .c(n859) );
	inv_0 U2799 ( .x(n861), .a(n816) );
	inv_8 U28 ( .x(net151622), .a(___cell__39620_net143983) );
	nor2i_3 U280 ( .x(n1039), .a(n855), .b(n1040) );
	aoi222_1 U2800 ( .x(n2936), .a(n1191), .b(n2859), .c(n650), .d(n2899),
		.e(n1221), .f(n2902) );
	aoi22_1 U2801 ( .x(n2901), .a(n1221), .b(n2863), .c(n1191), .d(n2902) );
	or3i_5 U2802 ( .x(n2295), .a(n2296), .b(n2293), .c(n864) );
	ao21_3 U2803 ( .x(n864), .a(n1085), .b(n2290), .c(n2291) );
	inv_12 U2804 ( .x(n3629), .a(n3628) );
	oai21_1 U2805 ( .x(n866), .a(n1587), .b(n889), .c(n3786) );
	oai21_1 U2806 ( .x(n867), .a(n1587), .b(n546), .c(n3786) );
	inv_2 U2807 ( .x(n3788), .a(n3787) );
	mux2_4 U2808 ( .x(n868), .d0(n3358), .sl(n816), .d1(n3313) );
	nand2i_2 U2809 ( .x(n3920), .a(n1632), .b(n827) );
	nand2i_0 U281 ( .x(n3616), .a(n1578), .b(n896) );
	and4i_2 U2810 ( .x(n2117), .a(n2116), .b(n2118), .c(n2119), .d(n2120) );
	oa211_5 U2811 ( .x(n869), .a(n844), .b(n4005), .c(n2632), .d(n3838) );
	inv_5 U2812 ( .x(n2107), .a(n870) );
	inv_14 U2813 ( .x(n872), .a(n874) );
	aoi221_1 U2814 ( .x(n2793), .a(n842), .b(n502), .c(___cell__39620_net143722),
		.d(n2798), .e(n1266) );
	aoi21_3 U2815 ( .x(n2675), .a(n2676), .b(n2677), .c(n2634) );
	oa22_4 U2816 ( .x(n2267), .a(n1730), .b(n877), .c(n1175), .d(n876) );
	inv_0 U2817 ( .x(n876), .a(n904) );
	inv_0 U2818 ( .x(n877), .a(n919) );
	nand2i_3 U2819 ( .x(n1730), .a(n1565), .b(n1689) );
	nand2_2 U282 ( .x(n3556), .a(n1040), .b(n3616) );
	inv_16 U2820 ( .x(n881), .a(n1643) );
	nand2i_2 U2821 ( .x(n3969), .a(n1634), .b(n525) );
	buf_1 U2822 ( .x(n919), .a(n931) );
	oaoi211_1 U2823 ( .x(n2606), .a(n2607), .b(n1700), .c(n541), .d(n2604) );
	oai21_1 U2824 ( .x(n2288), .a(n3737), .b(n1700), .c(reg_out_A[31]) );
	oai21_1 U2825 ( .x(n2486), .a(n3792), .b(n1700), .c(n537) );
	aoi21_1 U2826 ( .x(n3144), .a(n901), .b(n1700), .c(n1404) );
	aoi222_1 U2827 ( .x(n3053), .a(n1204), .b(n3056), .c(n644), .d(n1700),
		.e(ALU_result[14]), .f(n3057) );
	aoi21_1 U2828 ( .x(n2799), .a(n749), .b(n1700), .c(n1269) );
	oai21_1 U2829 ( .x(n2656), .a(n3841), .b(n1700), .c(n636) );
	inv_2 U283 ( .x(n3492), .a(n3647) );
	oai21_1 U2830 ( .x(n2530), .a(n3805), .b(n1700), .c(n540) );
	aoi21_1 U2831 ( .x(n3014), .a(n609), .b(n1700), .c(n1347) );
	aoi21_1 U2832 ( .x(n2978), .a(n893), .b(n1700), .c(n1328) );
	oai21_1 U2833 ( .x(n2697), .a(n3848), .b(n1700), .c(n686) );
	aoi21_1 U2834 ( .x(n2254), .a(n834), .b(n1700), .c(n1145) );
	aoi21_1 U2835 ( .x(n2105), .a(n852), .b(n1700), .c(n1107) );
	nand2i_1 U2836 ( .x(n2032), .a(n1529), .b(n1700) );
	aoi21_1 U2837 ( .x(n2063), .a(n914), .b(n1700), .c(n1086) );
	aoi21_1 U2838 ( .x(n2154), .a(n838), .b(n1700), .c(n1118) );
	inv_16 U2839 ( .x(n888), .a(n1652) );
	buf_3 U284 ( .x(n687), .a(reg_out_A[22]) );
	inv_16 U2840 ( .x(n891), .a(n1602) );
	buf_16 U2841 ( .x(n922), .a(n937) );
	exnor2_1 U2842 ( .x(n1492), .a(n628), .b(Imm[21]) );
	nand2_0 U2843 ( .x(n2720), .a(Imm[21]), .b(n628) );
	inv_0 U2844 ( .x(___cell__39620_net144765), .a(Imm[21]) );
	inv_16 U2845 ( .x(n894), .a(n1579) );
	nand2i_4 U2846 ( .x(n1652), .a(n891), .b(n531) );
	nand2_0 U2847 ( .x(___cell__39620_net146131), .a(n631), .b(n893) );
	exnor2_1 U2848 ( .x(n1504), .a(n893), .b(n631) );
	inv_0 U2849 ( .x(n898), .a(n904) );
	nand2i_2 U285 ( .x(n2605), .a(n1485), .b(n2139) );
	exnor2_1 U2850 ( .x(n1507), .a(net156363), .b(n644) );
	nand2_0 U2851 ( .x(n3023), .a(net156363), .b(n644) );
	inv_14 U2852 ( .x(n917), .a(n916) );
	inv_16 U2853 ( .x(n904), .a(n903) );
	nand2i_2 U2854 ( .x(n3354), .a(n1585), .b(n839) );
	nand2i_2 U2855 ( .x(n3555), .a(n1648), .b(n839) );
	nand2i_2 U2856 ( .x(n3564), .a(n862), .b(n839) );
	nand2i_2 U2857 ( .x(n3309), .a(n1561), .b(n839) );
	nand2i_2 U2858 ( .x(n3348), .a(n1563), .b(n839) );
	nand2i_2 U2859 ( .x(n3500), .a(n1577), .b(n839) );
	oai221_1 U286 ( .x(n3523), .a(n1302), .b(n1043), .c(n3524), .d(n4007),
		.e(n1806) );
	nand2i_2 U2860 ( .x(n3405), .a(n748), .b(n839) );
	nand2i_2 U2861 ( .x(n3338), .a(n1579), .b(n839) );
	nand2i_2 U2862 ( .x(n3474), .a(n1570), .b(n839) );
	nand2i_2 U2863 ( .x(n3353), .a(n1571), .b(n839) );
	nand2i_2 U2864 ( .x(n3320), .a(n1572), .b(n839) );
	nand2i_2 U2865 ( .x(n3329), .a(n1586), .b(n839) );
	nand2i_2 U2866 ( .x(n3495), .a(n1583), .b(n839) );
	nand2i_2 U2867 ( .x(n3491), .a(n1584), .b(n839) );
	inv_16 U2868 ( .x(n910), .a(n909) );
	exnor2_1 U2869 ( .x(n1510), .a(reg_out_B[13]), .b(n919) );
	and2_3 U287 ( .x(n733), .a(IR_opcode_field[3]), .b(IR_opcode_field[2]) );
	nand2_1 U2870 ( .x(n2260), .a(n3573), .b(n919) );
	inv_2 U2871 ( .x(n1563), .a(n930) );
	buf_1 U2872 ( .x(n920), .a(n937) );
	inv_16 U2873 ( .x(n914), .a(n913) );
	inv_0 U2874 ( .x(n945), .a(reg_dst) );
	aoai211_3 U2875 ( .x(n4116), .a(n946), .b(n947), .c(reg_dst), .d(N3304) );
	exnor2_1 U2876 ( .x(n1509), .a(n629), .b(n919) );
	nor2i_0 U2877 ( .x(n3060), .a(n629), .b(n1563) );
	inv_0 U2878 ( .x(n1375), .a(n629) );
	exnor2_1 U2879 ( .x(n1511), .a(n682), .b(n894) );
	nand3_0 U288 ( .x(___cell__39620_net143836), .a(n733), .b(n1520), .c(___cell__39620_net144355) );
	nor2i_0 U2880 ( .x(n1377), .a(n682), .b(n1579) );
	inv_6 U2881 ( .x(n916), .a(n4015) );
	inv_2 U2882 ( .x(n1037), .a(counter[1]) );
	inv_10 U2883 ( .x(n937), .a(n935) );
	mux2i_5 U2884 ( .x(n3172), .d0(n3531), .sl(net149120), .d1(n3446) );
	inv_10 U2885 ( .x(n3531), .a(n3530) );
	nand2_0 U2886 ( .x(n2112), .a(n838), .b(n642) );
	inv_0 U2887 ( .x(___cell__39620_net143735), .a(n642) );
	exnor2_1 U2888 ( .x(n1463), .a(n642), .b(n922) );
	inv_0 U2889 ( .x(n1208), .a(n818) );
	inv_5 U289 ( .x(n2079), .a(n1682) );
	nor2i_0 U2890 ( .x(n1406), .a(n818), .b(n1572) );
	exnor2_1 U2891 ( .x(n1516), .a(n818), .b(n908) );
	nand2i_0 U2892 ( .x(n1610), .a(IR_opcode_field[3]), .b(IR_opcode_field[2]) );
	oai21_1 U2895 ( .x(n3238), .a(n1166), .b(n546), .c(n3239) );
	oai21_1 U2896 ( .x(n3787), .a(n1587), .b(n889), .c(n3786) );
	nand3i_3 U2897 ( .x(n4050), .a(n948), .b(n949), .c(n950) );
	oai211_4 U2898 ( .x(n4051), .a(n951), .b(___cell__39620_net147731), .c(n952),
		.d(n953) );
	oai211_3 U2899 ( .x(n4054), .a(n954), .b(___cell__39620_net147731), .c(n955),
		.d(n956) );
	inv_8 U29 ( .x(n684), .a(n683) );
	inv_4 U290 ( .x(n3202), .a(n695) );
	nand2_2 U2900 ( .x(n4065), .a(n972), .b(n973) );
	nand4_1 U2901 ( .x(n4074), .a(n983), .b(n984), .c(n985), .d(n986) );
	nand3i_3 U2902 ( .x(n4079), .a(n554), .b(n994), .c(n995) );
	nand2i_4 U2903 ( .x(n4073), .a(n1015), .b(n1016) );
	nand2_2 U2904 ( .x(n4066), .a(n1026), .b(n1027) );
	oai211_4 U2905 ( .x(n4064), .a(n1028), .b(___cell__39620_net143287), .c(n1029),
		.d(n1030) );
	oai211_3 U2906 ( .x(n4062), .a(n1031), .b(___cell__39620_net143287), .c(n1032),
		.d(n1033) );
	nor2i_5 U2907 ( .x(n1053), .a(n1054), .b(n1055) );
	nor2i_5 U2908 ( .x(n1068), .a(n1069), .b(n4004) );
	nor2_6 U2909 ( .x(n1097), .a(n947), .b(n1098) );
	and4i_4 U2910 ( .x(n957), .a(n1103), .b(n1100), .c(n1101), .d(n1102) );
	nor2i_5 U2911 ( .x(n1108), .a(n922), .b(n1089) );
	nor2i_5 U2912 ( .x(n1135), .a(n1136), .b(n4007) );
	and4i_4 U2913 ( .x(n1001), .a(n1141), .b(n1138), .c(n1139), .d(n1140) );
	and4i_4 U2914 ( .x(n1004), .a(n1173), .b(n1170), .c(n1171), .d(n1172) );
	nor2_6 U2915 ( .x(n1180), .a(n679), .b(n4037) );
	nor2i_5 U2916 ( .x(n1183), .a(N1959), .b(n1184) );
	nor2i_5 U2917 ( .x(n1187), .a(n590), .b(n1120) );
	nor2i_5 U2918 ( .x(n1193), .a(n541), .b(n1120) );
	nor2i_5 U2919 ( .x(n1194), .a(n541), .b(n1122) );
	oai22_1 U292 ( .x(n2564), .a(n1578), .b(n695), .c(n2565), .d(n1682) );
	nor2i_5 U2920 ( .x(n1195), .a(N1957), .b(n1184) );
	and4i_4 U2921 ( .x(n987), .a(n1202), .b(n1199), .c(n1200), .d(n1201) );
	aoi21_3 U2922 ( .x(n1015), .a(n1231), .b(n1232), .c(___cell__39620_net147731) );
	nor2i_5 U2923 ( .x(n1251), .a(N1984), .b(___cell__39620_net143845) );
	nor2i_5 U2924 ( .x(n1293), .a(N2015), .b(n1169) );
	nor2_6 U2925 ( .x(n1305), .a(n947), .b(n1306) );
	nor2i_5 U2926 ( .x(n1307), .a(n1308), .b(n1166) );
	nor2i_5 U2927 ( .x(n1338), .a(n1339), .b(n1055) );
	and4i_4 U2928 ( .x(n969), .a(n1355), .b(n1352), .c(n1353), .d(n1354) );
	and4i_4 U2929 ( .x(n1031), .a(n1368), .b(n1365), .c(n1366), .d(n1367) );
	nand2i_5 U293 ( .x(n4012), .a(n1556), .b(reg_out_B[3]) );
	and4i_4 U2930 ( .x(n966), .a(n1386), .b(n1383), .c(n1384), .d(n1385) );
	nor2i_5 U2931 ( .x(n1433), .a(n1434), .b(___cell__39620_net143653) );
	nand2i_4 U2932 ( .x(n1541), .a(n1534), .b(n1542) );
	nand2i_4 U2933 ( .x(n1070), .a(reg_out_B[3]), .b(n815) );
	inv_6 U2935 ( .x(n1572), .a(n908) );
	nand3i_5 U2936 ( .x(n1169), .a(___cell__39620_net143653), .b(n810), .c(n1520) );
	nand2i_4 U2937 ( .x(___cell__39620_net144340), .a(n1610), .b(n4137) );
	or3i_5 U2938 ( .x(___cell__39620_net144343), .a(___cell__39620_net144344),
		.b(net152465), .c(___cell__39620_net143653) );
	nand2i_4 U2939 ( .x(n1620), .a(n1621), .b(n676) );
	exnor2_1 U294 ( .x(n1484), .a(n590), .b(reg_out_B[25]) );
	nand2i_4 U2940 ( .x(n1627), .a(n1628), .b(n1543) );
	or2_8 U2942 ( .x(n1636), .a(n816), .b(n815) );
	inv_6 U2943 ( .x(n1098), .a(N1870) );
	inv_6 U2944 ( .x(n1736), .a(N1893) );
	oai21_5 U2945 ( .x(n1740), .a(n1642), .b(n1654), .c(n1741) );
	inv_6 U2946 ( .x(n1775), .a(N1658) );
	inv_6 U2947 ( .x(n1778), .a(N1823) );
	inv_6 U2948 ( .x(n1780), .a(N1856) );
	inv_6 U2949 ( .x(n1820), .a(N1752) );
	nand2_2 U295 ( .x(n2283), .a(n3499), .b(n3500) );
	oai21_4 U2950 ( .x(n1939), .a(n1531), .b(n1940), .c(n1447) );
	mux2i_3 U2951 ( .x(n4080), .d0(n4047), .sl(N3304), .d1(n1941) );
	mux2i_3 U2952 ( .x(n4048), .d0(n4046), .sl(N3304), .d1(n1942) );
	inv_6 U2953 ( .x(n1434), .a(N3024) );
	mux2i_3 U2954 ( .x(n1943), .d0(N3024), .sl(IR_opcode_field[0]), .d1(N3029) );
	mux2i_3 U2955 ( .x(n1944), .d0(n1945), .sl(IR_opcode_field[1]), .d1(n1946) );
	inv_6 U2956 ( .x(n1947), .a(N1392) );
	mux2i_3 U2957 ( .x(n1948), .d0(N1402), .sl(IR_function_field[0]), .d1(N1407) );
	nand2i_4 U2958 ( .x(___cell__39620_net144173), .a(IR_opcode_field[1]),
		.b(___cell__39620_net145037) );
	nor2_5 U2959 ( .x(n1549), .a(n1956), .b(n1957) );
	inv_2 U296 ( .x(n2183), .a(n1713) );
	aoi22_3 U2960 ( .x(n1963), .a(n1964), .b(n1965), .c(n1330), .d(n1966) );
	nor2i_5 U2961 ( .x(n1575), .a(n1451), .b(___cell__39620_net144175) );
	nor2_6 U2962 ( .x(n1581), .a(___cell__39620_net144175), .b(n1451) );
	aoi22_3 U2963 ( .x(n1975), .a(n1964), .b(n1976), .c(n1330), .d(n1977) );
	nand4_1 U2964 ( .x(n1059), .a(n1989), .b(n1990), .c(n1986), .d(n1991) );
	oai22_3 U2965 ( .x(n2010), .a(n2011), .b(n1574), .c(n2012), .d(n1566) );
	and4i_4 U2966 ( .x(n962), .a(n2010), .b(n2013), .c(n2015), .d(n2016) );
	and4i_4 U2967 ( .x(n961), .a(n2020), .b(n2017), .c(n2018), .d(n2019) );
	nand4_1 U2968 ( .x(n1081), .a(n2040), .b(n2041), .c(n2039), .d(n2042) );
	nand2_2 U297 ( .x(n2284), .a(n3404), .b(n3405) );
	oai211_4 U2970 ( .x(n2056), .a(n580), .b(n621), .c(n2060), .d(n2061) );
	aoi211_5 U2971 ( .x(n2058), .a(n1204), .b(n2064), .c(n1084), .d(n2062) );
	nand2i_4 U2972 ( .x(n1676), .a(net149167), .b(net151904) );
	aoi211_4 U2973 ( .x(n2078), .a(n2079), .b(n2080), .c(n1088), .d(n1090) );
	nand4_1 U2974 ( .x(n2097), .a(n2100), .b(n2101), .c(n2102), .d(n2098) );
	oai21_5 U2975 ( .x(n2111), .a(n881), .b(n1644), .c(n2110) );
	ao221_4 U2976 ( .x(n2121), .a(n662), .b(n1993), .c(n1318), .d(n2043), .e(n1112) );
	oai211_3 U2977 ( .x(n2143), .a(n2012), .b(n1186), .c(n2144), .d(n2145) );
	nor2i_5 U2978 ( .x(n2162), .a(n2163), .b(n1982) );
	and4i_4 U2979 ( .x(n1126), .a(n2171), .b(n2173), .c(n2174), .d(n2175) );
	and2_3 U298 ( .x(n507), .a(n3540), .b(n522) );
	aoi21_3 U2980 ( .x(n2180), .a(n1391), .b(n2181), .c(n1119) );
	and3i_3 U2981 ( .x(n955), .a(n2198), .b(n2200), .c(n2201) );
	and3i_3 U2982 ( .x(n2202), .a(n2205), .b(n2203), .c(n2204) );
	aoi21_3 U2983 ( .x(n2220), .a(n1318), .b(n2168), .c(n1137) );
	nand4_1 U2984 ( .x(n1141), .a(n2219), .b(n2217), .c(n2221), .d(n2220) );
	aoi21_3 U2985 ( .x(n2229), .a(n1066), .b(n2045), .c(n1133) );
	and3i_3 U2986 ( .x(n1002), .a(n2242), .b(n2244), .c(n2245) );
	nand4_1 U2987 ( .x(n2248), .a(n2249), .b(n2250), .c(n2251), .d(n2252) );
	nor2i_3 U2988 ( .x(n2245), .a(n2246), .b(n2253) );
	nand4_1 U2989 ( .x(n2253), .a(n2255), .b(n2256), .c(n2254), .d(n2257) );
	inv_14 U299 ( .x(n1689), .a(n1633) );
	nor2i_5 U2990 ( .x(___cell__39620_net145450), .a(n1683), .b(n1626) );
	aoi22_3 U2991 ( .x(n2301), .a(___cell__39620_net144517), .b(n2302), .c(n1391),
		.d(n2303) );
	nand4_1 U2992 ( .x(n2325), .a(___cell__39620_net145470), .b(n2326), .c(n2323),
		.d(n2317) );
	aoi21_3 U2993 ( .x(n2342), .a(n1177), .b(n1977), .c(n2067) );
	and4i_5 U2994 ( .x(n1170), .a(n1164), .b(n2350), .c(n2351), .d(n2346) );
	oai22_3 U2995 ( .x(n2358), .a(n2359), .b(n1588), .c(n2360), .d(n1574) );
	and4i_4 U2996 ( .x(n1006), .a(n2358), .b(n2361), .c(n2362), .d(n2363) );
	aoi21_3 U2998 ( .x(n2437), .a(n1066), .b(n2303), .c(n1187) );
	nand4_1 U2999 ( .x(n2443), .a(n2446), .b(n2447), .c(n2448), .d(n2449) );
	buf_10 U3 ( .x(net149121), .a(net149107) );
	inv_2 U30 ( .x(net156024), .a(Imm[17]) );
	nand4_1 U3000 ( .x(n2450), .a(n2453), .b(n2452), .c(n2451), .d(n2454) );
	nor3_4 U3001 ( .x(n1008), .a(n2450), .b(n2442), .c(n2438) );
	nand2_5 U3002 ( .x(n2459), .a(n1267), .b(___cell__39620_net144345) );
	oai221_3 U3003 ( .x(n2463), .a(___cell__39620_net143872), .b(n1764), .c(___cell__39620_net143660),
		.d(n1765), .e(n2464) );
	oai211_3 U3004 ( .x(n2466), .a(n553), .b(n1055), .c(n2467), .d(n2468) );
	nand4_1 U3005 ( .x(n1202), .a(n2469), .b(n2470), .c(n2471), .d(n2472) );
	aoi21_3 U3006 ( .x(n2480), .a(n1066), .b(n2375), .c(n1193) );
	nand4i_4 U3007 ( .x(n2497), .a(n1203), .b(n2498), .c(n2500), .d(n2501) );
	and4i_4 U3008 ( .x(n2504), .a(n2507), .b(n2505), .c(n2506), .d(n2503) );
	aoi22_3 U3009 ( .x(n2519), .a(n2079), .b(n2262), .c(n1391), .d(n2520) );
	inv_5 U301 ( .x(n1219), .a(reg_out_A[25]) );
	aoi21_3 U3010 ( .x(n2522), .a(___cell__39620_net144517), .b(n2303), .c(n2521) );
	and4i_4 U3011 ( .x(n1012), .a(n2527), .b(n2533), .c(n2534), .d(n2531) );
	and4i_4 U3012 ( .x(n1011), .a(n2538), .b(n2535), .c(n2536), .d(n2537) );
	nor2i_5 U3013 ( .x(n2535), .a(n2539), .b(n1210) );
	and4i_4 U3014 ( .x(n2577), .a(n2575), .b(n2567), .c(n2569), .d(n2573) );
	and3i_3 U3015 ( .x(n983), .a(n2579), .b(n2578), .c(n2577) );
	nor3i_5 U3016 ( .x(n2578), .a(n2585), .b(n1223), .c(n1225) );
	nand2_5 U3017 ( .x(n2589), .a(n2590), .b(n2591) );
	nand3i_3 U3018 ( .x(n2598), .a(n1229), .b(n2601), .c(n2599) );
	oai211_3 U3019 ( .x(n2610), .a(n2611), .b(n1186), .c(n2606), .d(n2608) );
	nand2_6 U302 ( .x(n1091), .a(n1686), .b(n1683) );
	aoi21_3 U3020 ( .x(n2612), .a(n1191), .b(n2532), .c(n2613) );
	and3i_3 U3021 ( .x(n2616), .a(n2619), .b(n2621), .c(n2622) );
	aoi21_3 U3022 ( .x(n2623), .a(___cell__39620_net143722), .b(n2624), .c(n1233) );
	nand4_1 U3023 ( .x(n2636), .a(n2637), .b(n2638), .c(n2639), .d(n2635) );
	oai211_3 U3024 ( .x(n2643), .a(n869), .b(n1166), .c(n2644), .d(n2645) );
	and3i_4 U3025 ( .x(n1238), .a(n2643), .b(n2646), .c(n2647) );
	aoi22_4 U3026 ( .x(n2648), .a(n1683), .b(n2375), .c(___cell__39620_net144517),
		.d(n2649) );
	aoi21_6 U3027 ( .x(n2682), .a(n2674), .b(___cell__39620_net147791), .c(n1241) );
	nand4_1 U3028 ( .x(n1247), .a(n2685), .b(n2686), .c(n2687), .d(n2688) );
	oai211_3 U3029 ( .x(n2695), .a(n2696), .b(n1566), .c(n2692), .d(n2697) );
	oai22_1 U303 ( .x(n2521), .a(n1529), .b(n1091), .c(n1219), .d(n695) );
	and4i_4 U3030 ( .x(n2700), .a(n2695), .b(n2701), .c(n2702), .d(n2698) );
	nand4_1 U3031 ( .x(n2705), .a(n2715), .b(n2716), .c(n2717), .d(n2712) );
	aoi22_4 U3032 ( .x(n2740), .a(n2139), .b(n2741), .c(n2193), .d(n2742) );
	oai22_3 U3033 ( .x(n2745), .a(n2696), .b(n1574), .c(n2746), .d(n1566) );
	oai22_3 U3034 ( .x(n2748), .a(n1143), .b(n1816), .c(n2655), .d(n1588) );
	and3i_3 U3035 ( .x(n2751), .a(n2753), .b(n2757), .c(n2758) );
	and4i_4 U3036 ( .x(n2768), .a(n2772), .b(n2769), .c(n2770), .d(n2771) );
	oai22_3 U3037 ( .x(n2791), .a(___cell__39620_net143693), .b(___cell__39620_net144781),
		.c(n2696), .d(n1588) );
	nor3_4 U3038 ( .x(n2792), .a(n2791), .b(n2788), .c(n2789) );
	nand4_1 U3039 ( .x(n2795), .a(n2799), .b(n2800), .c(n2801), .d(n2796) );
	inv_5 U304 ( .x(n1528), .a(n1525) );
	aoi21_6 U3040 ( .x(n2810), .a(n1177), .b(n1969), .c(n1836) );
	nand4_1 U3041 ( .x(n1277), .a(n2813), .b(n2815), .c(n2816), .d(n2814) );
	aoi221_4 U3042 ( .x(n2817), .a(n1095), .b(n1423), .c(n1197), .d(n1165),
		.e(n1273) );
	nand4_3 U3043 ( .x(n1276), .a(n2817), .b(n2818), .c(n2819), .d(n2820) );
	oai211_4 U3044 ( .x(n2821), .a(n2822), .b(n1626), .c(n2823), .d(n2824) );
	nand4_3 U3045 ( .x(n2830), .a(n2831), .b(n2832), .c(n2828), .d(n2833) );
	nor3_4 U3046 ( .x(n952), .a(n2821), .b(n2830), .c(n2825) );
	and3i_3 U3048 ( .x(n2896), .a(n2893), .b(n2891), .c(n2897) );
	and3i_3 U3049 ( .x(n2903), .a(n2898), .b(n2901), .c(n2904) );
	nand2i_0 U305 ( .x(n2460), .a(reg_out_B[4]), .b(n1964) );
	and4i_4 U3050 ( .x(n2918), .a(n1317), .b(n2917), .c(n2919), .d(n2914) );
	nand3i_3 U3051 ( .x(n2937), .a(n2931), .b(n2928), .c(n2936) );
	oai22_3 U3052 ( .x(n2942), .a(n2943), .b(n1658), .c(n2944), .d(n784) );
	ao21_4 U3053 ( .x(n2941), .a(n1085), .b(n2910), .c(n2945) );
	ao21_4 U3054 ( .x(n2961), .a(n1221), .b(n2859), .c(n2958) );
	nand4_1 U3055 ( .x(n2966), .a(n2967), .b(n2968), .c(n2965), .d(n2969) );
	and3i_3 U3056 ( .x(n973), .a(n2966), .b(n2962), .c(n2970) );
	nand2_5 U3057 ( .x(n2971), .a(n2972), .b(n2973) );
	and4i_4 U3058 ( .x(n2968), .a(n2971), .b(n2974), .c(n2975), .d(n2976) );
	and3i_4 U3059 ( .x(n2967), .a(n2977), .b(n2978), .c(n2979) );
	nor2i_3 U306 ( .x(n2458), .a(___cell__39620_net144331), .b(n1072) );
	and4i_5 U3060 ( .x(n1342), .a(n1338), .b(n2982), .c(n2983), .d(n2984) );
	nand3_3 U3061 ( .x(n3005), .a(n3002), .b(n2999), .c(n3003) );
	and4i_4 U3062 ( .x(n3015), .a(n3018), .b(n3016), .c(n3017), .d(n3014) );
	nand4_1 U3063 ( .x(n1355), .a(n3029), .b(n3030), .c(n3028), .d(n3031) );
	nand4i_4 U3064 ( .x(n3045), .a(n3037), .b(n3039), .c(n3044), .d(n3046) );
	nand4_1 U3065 ( .x(n3048), .a(n3052), .b(n3053), .c(n3049), .d(n3050) );
	nand4_1 U3066 ( .x(n1368), .a(n3064), .b(n3065), .c(n3066), .d(n3067) );
	aoi221_4 U3067 ( .x(n3074), .a(___cell__39620_net143864), .b(n3075), .c(___cell__39620_net143722),
		.d(n3076), .e(n1372) );
	aoi221_4 U3068 ( .x(n3077), .a(n650), .b(n3041), .c(n649), .d(n3078), .e(n3079) );
	nor3_4 U3069 ( .x(n3082), .a(n3083), .b(n3084), .c(n3085) );
	nand2i_2 U307 ( .x(___cell__39620_net144200), .a(n1533), .b(IR_opcode_field[1]) );
	nand4i_4 U3071 ( .x(n3105), .a(n3099), .b(n3101), .c(n3104), .d(n3106) );
	nand4_1 U3072 ( .x(n1402), .a(n3123), .b(n3124), .c(n3122), .d(n3125) );
	and4i_4 U3073 ( .x(n1410), .a(n3149), .b(n3151), .c(n3148), .d(n3152) );
	oai22_3 U3074 ( .x(n3160), .a(n3130), .b(n1574), .c(n2011), .d(n1566) );
	ao21_4 U3075 ( .x(n3185), .a(n1066), .b(n3186), .c(n3182) );
	and4i_5 U3076 ( .x(n3192), .a(n1422), .b(n3193), .c(n3194), .d(n3191) );
	oai211_3 U3077 ( .x(n3203), .a(n3204), .b(n3180), .c(n3205), .d(n3206) );
	oai211_3 U3078 ( .x(n3208), .a(n2360), .b(n1186), .c(n3209), .d(n3210) );
	nor3_4 U3079 ( .x(n949), .a(n3203), .b(n3208), .c(n3207) );
	nand2_2 U308 ( .x(n3315), .a(n1040), .b(n3595) );
	nand4_1 U3080 ( .x(n3220), .a(n1514), .b(n1511), .c(n1516), .d(n1517) );
	nand4_1 U3081 ( .x(n3223), .a(n1497), .b(n1495), .c(n1501), .d(n1499) );
	nand4_1 U3082 ( .x(n3224), .a(n1490), .b(n1488), .c(n1494), .d(n1492) );
	nand4_1 U3083 ( .x(n3226), .a(n1481), .b(n1479), .c(n1486), .d(n1483) );
	nand4_1 U3084 ( .x(n3227), .a(n1473), .b(n1471), .c(n1477), .d(n1475) );
	nand4_1 U3085 ( .x(n3229), .a(n1465), .b(n1463), .c(n1469), .d(n1467) );
	nor3i_5 U3086 ( .x(n3246), .a(n3247), .b(n3242), .c(n1435) );
	nand3_3 U3087 ( .x(n1441), .a(n3246), .b(n3244), .c(n3248) );
	nand4_1 U3088 ( .x(n3261), .a(n1498), .b(n1496), .c(n1502), .d(n1500) );
	nand4_1 U3089 ( .x(n3262), .a(n1489), .b(n1487), .c(n1493), .d(n1491) );
	inv_2 U309 ( .x(n3595), .a(n651) );
	nand4_1 U3090 ( .x(n3264), .a(n1482), .b(n1480), .c(n1485), .d(n1484) );
	nand4_1 U3091 ( .x(n3272), .a(n1466), .b(n1464), .c(n1470), .d(n1468) );
	nand4_1 U3092 ( .x(n3273), .a(n1461), .b(n1459), .c(n3274), .d(n1457) );
	aoi211_4 U3093 ( .x(n3282), .a(n3283), .b(n2004), .c(n1449), .d(n3284) );
	nand2_5 U3094 ( .x(n3291), .a(n3292), .b(n3293) );
	ao211_5 U3095 ( .x(n1966), .a(reg_out_B[4]), .b(n3311), .c(n897), .d(n2067) );
	oai22_5 U3096 ( .x(n3312), .a(n915), .b(n1654), .c(n1642), .d(n1655) );
	ao211_5 U3097 ( .x(n1969), .a(reg_out_B[4]), .b(n3315), .c(n3316), .d(n2067) );
	inv_5 U3098 ( .x(n3324), .a(n3321) );
	ao211_5 U3099 ( .x(n1977), .a(reg_out_B[4]), .b(n3325), .c(n3326), .d(n2067) );
	inv_2 U31 ( .x(n639), .a(n638) );
	nand2_2 U310 ( .x(n3351), .a(n1040), .b(n3596) );
	ao211_5 U3100 ( .x(n1069), .a(reg_out_B[4]), .b(n3332), .c(n3333), .d(n2067) );
	ao211_5 U3101 ( .x(n1965), .a(reg_out_B[4]), .b(n3343), .c(n3344), .d(n2067) );
	nand2i_4 U3102 ( .x(n1976), .a(n1973), .b(n3354) );
	nand2_5 U3103 ( .x(n2992), .a(n3370), .b(n3371) );
	oai22_5 U3104 ( .x(n2568), .a(n1573), .b(n1642), .c(___cell__39620_net144257),
		.d(n915) );
	oai22_3 U3105 ( .x(n2306), .a(n509), .b(n536), .c(n1585), .d(n1629) );
	oai22_3 U3106 ( .x(n2373), .a(n3409), .b(n536), .c(n1571), .d(n1629) );
	oai211_4 U3107 ( .x(n3422), .a(n3423), .b(n1560), .c(n3424), .d(n3425) );
	oai22_3 U3108 ( .x(n2738), .a(n507), .b(reg_out_B[3]), .c(n1572), .d(n822) );
	oai22_3 U3109 ( .x(n2477), .a(n3406), .b(n536), .c(n1579), .d(n1629) );
	nand2i_2 U311 ( .x(n1157), .a(N69), .b(n1552) );
	oai22_5 U3111 ( .x(n2375), .a(n1571), .b(n871), .c(n3454), .d(n4125) );
	oai22_5 U3112 ( .x(n3457), .a(n1561), .b(n872), .c(net149167), .d(n3341) );
	oai22_3 U3113 ( .x(n3458), .a(n1529), .b(n872), .c(n3459), .d(n4125) );
	nand2i_4 U3114 ( .x(n3464), .a(n3465), .b(n3466) );
	nand2i_4 U3115 ( .x(n3467), .a(n3468), .b(n3469) );
	ao211_5 U3116 ( .x(n1349), .a(net151904), .b(n3477), .c(n547), .d(n1982) );
	ao211_5 U3117 ( .x(n1047), .a(net151904), .b(n3478), .c(n3322), .d(n1982) );
	ao211_5 U3118 ( .x(n1049), .a(net151904), .b(n3479), .c(n3468), .d(n1982) );
	ao211_5 U3119 ( .x(n1045), .a(net151904), .b(n3480), .c(n622), .d(n1982) );
	nor2i_0 U312 ( .x(n1156), .a(n855), .b(n1157) );
	ao211_5 U3120 ( .x(n1361), .a(net151904), .b(n3482), .c(n3471), .d(n1982) );
	nand2i_4 U3121 ( .x(n3496), .a(n3497), .b(n3498) );
	oai221_3 U3122 ( .x(n2167), .a(n3509), .b(n1607), .c(n891), .d(n3510),
		.e(n3511) );
	ao221_5 U3123 ( .x(n2165), .a(n1289), .b(n3537), .c(n3186), .d(n1602),
		.e(n1123) );
	ao221_5 U3124 ( .x(n2218), .a(n1289), .b(n3538), .c(n3539), .d(n1602),
		.e(n1135) );
	nand2i_4 U3125 ( .x(n3541), .a(n3542), .b(n3543) );
	oai22_5 U3126 ( .x(n3544), .a(n1572), .b(n880), .c(n822), .d(n1646) );
	ao211_5 U3127 ( .x(n3278), .a(reg_out_B[4]), .b(n3556), .c(n2067), .d(n3557) );
	ao211_5 U3128 ( .x(n1136), .a(net151904), .b(n3559), .c(n1982), .d(n3558) );
	nand2_5 U3129 ( .x(n3560), .a(n3561), .b(n3562) );
	nand2_2 U313 ( .x(n3783), .a(n3325), .b(n855) );
	oai22_5 U3130 ( .x(n2179), .a(n557), .b(n836), .c(n3489), .d(n4125) );
	nand2i_4 U3131 ( .x(n3570), .a(n1562), .b(n1728) );
	inv_5 U3132 ( .x(n3322), .a(n3574) );
	inv_5 U3133 ( .x(n3471), .a(n3578) );
	inv_5 U3134 ( .x(n3465), .a(n3588) );
	inv_5 U3135 ( .x(n3468), .a(n3589) );
	inv_5 U3136 ( .x(n3605), .a(n3495) );
	nand2i_4 U3138 ( .x(n1606), .a(net151904), .b(n1982) );
	inv_5 U3139 ( .x(n3389), .a(n3637) );
	nand2_2 U314 ( .x(n3332), .a(n1040), .b(n3615) );
	inv_5 U3140 ( .x(n3542), .a(n3657) );
	nand2i_4 U3142 ( .x(n3682), .a(n1655), .b(n883) );
	oai211_3 U3143 ( .x(n3683), .a(n1331), .b(n1546), .c(n2065), .d(n3682) );
	nand2_2 U3144 ( .x(n2100), .a(n2024), .b(n3669) );
	nand2i_4 U3146 ( .x(n3695), .a(n2114), .b(n3694) );
	nand4_1 U3147 ( .x(n999), .a(n2117), .b(n2122), .c(n3697), .d(n3696) );
	nand2i_4 U3148 ( .x(n2151), .a(n1626), .b(n3681) );
	nand2i_0 U315 ( .x(n3615), .a(n1580), .b(n896) );
	nand2i_4 U3150 ( .x(n3703), .a(n1561), .b(n2066) );
	nand2i_4 U3151 ( .x(n3704), .a(n1546), .b(n1965) );
	nand3_3 U3152 ( .x(n3176), .a(n3704), .b(n3703), .c(n2159) );
	inv_5 U3153 ( .x(n3436), .a(n3176) );
	oai22_5 U3154 ( .x(n3705), .a(n1660), .b(n1122), .c(n4001), .d(n1120) );
	nand3_3 U3155 ( .x(n3186), .a(n3707), .b(n3706), .c(n2162) );
	nand2i_4 U3156 ( .x(n2208), .a(n1626), .b(n3689) );
	nand3_3 U3157 ( .x(n3711), .a(n2229), .b(n3710), .c(n2228) );
	nand3_3 U3159 ( .x(n2371), .a(n2232), .b(n3712), .c(n2231) );
	nand2_2 U316 ( .x(n3802), .a(n3479), .b(___cell__39620_net144331) );
	nand2i_4 U3160 ( .x(n3713), .a(n748), .b(n2066) );
	nand2i_4 U3161 ( .x(n3714), .a(n1546), .b(n1069) );
	nand3_3 U3162 ( .x(n3715), .a(n3714), .b(n3713), .c(n2213) );
	inv_5 U3163 ( .x(n3430), .a(n3715) );
	nand2i_4 U3164 ( .x(n2250), .a(n1654), .b(___cell__39620_net145444) );
	nand4_3 U3166 ( .x(n3719), .a(n2282), .b(n3718), .c(n2281), .d(n3367) );
	oai21_4 U3167 ( .x(___cell__39620_net147270), .a(n3720), .b(n1451), .c(n2285) );
	nand2_5 U3168 ( .x(n2275), .a(n3573), .b(n894) );
	or3i_4 U3169 ( .x(___cell__39620_net145421), .a(___cell__39620_net147732),
		.b(n1169), .c(n1726) );
	nand2_2 U317 ( .x(n3481), .a(n665), .b(n3625) );
	or3i_4 U3170 ( .x(___cell__39620_net145425), .a(___cell__39620_net143326),
		.b(n1184), .c(n1727) );
	nand2_5 U3171 ( .x(n3392), .a(n1686), .b(n901) );
	aoai211_4 U3172 ( .x(___cell__39620_net145429), .a(n1545), .b(n3741), .c(n1158),
		.d(n619) );
	inv_5 U3173 ( .x(n3750), .a(n1740) );
	nand2i_4 U3174 ( .x(n3751), .a(n1560), .b(n3683) );
	nand3i_5 U3175 ( .x(n3752), .a(n1740), .b(n3751), .c(n2342) );
	nand4i_4 U3176 ( .x(n3755), .a(n1176), .b(n3750), .c(n2338), .d(n3416) );
	nand2i_4 U3177 ( .x(n2367), .a(n1657), .b(n3705) );
	inv_5 U3178 ( .x(n2439), .a(n3765) );
	nand3_3 U3179 ( .x(n2499), .a(n2431), .b(n3769), .c(n2430) );
	nand2_2 U318 ( .x(n3773), .a(n3481), .b(___cell__39620_net144331) );
	nand2i_4 U3180 ( .x(n3777), .a(n2460), .b(n1728) );
	nand2i_4 U3181 ( .x(n3781), .a(n4008), .b(n2279) );
	nand3_3 U3182 ( .x(n3785), .a(n2478), .b(n3784), .c(n2476) );
	nand3_3 U3183 ( .x(n3796), .a(n2519), .b(n3795), .c(n2522) );
	inv_5 U3184 ( .x(n1224), .a(n3796) );
	nand4_1 U3185 ( .x(n3800), .a(n2518), .b(n3797), .c(n3799), .d(n3798) );
	inv_5 U3186 ( .x(n1211), .a(n3800) );
	nand2i_4 U3187 ( .x(n3808), .a(n1626), .b(n867) );
	oai31_2 U3188 ( .x(n1014), .a(n2514), .b(n2508), .c(n1209), .d(___cell__39620_net147732) );
	nand4_1 U3189 ( .x(n3816), .a(n3814), .b(n3813), .c(n3815), .d(n2561) );
	nand2_2 U319 ( .x(n3482), .a(n665), .b(n3636) );
	inv_5 U3190 ( .x(n2670), .a(n2624) );
	oai211_3 U3191 ( .x(n3830), .a(n3553), .b(n1623), .c(n3829), .d(n2648) );
	inv_5 U3192 ( .x(n2667), .a(n3830) );
	oai211_3 U3193 ( .x(n2714), .a(n3460), .b(n4010), .c(n3843), .d(n2691) );
	oai211_3 U3194 ( .x(n2713), .a(n3403), .b(n1635), .c(n3844), .d(n2689) );
	nand2i_4 U3195 ( .x(n2701), .a(n1574), .b(n3837) );
	oai211_3 U3196 ( .x(n2803), .a(n3553), .b(n1625), .c(n3851), .d(n2739) );
	nand2i_4 U3197 ( .x(n3521), .a(n891), .b(n3033) );
	nand2_5 U3198 ( .x(n2827), .a(n2805), .b(n3864) );
	nand2i_4 U3199 ( .x(n2831), .a(n1186), .b(n2192) );
	inv_5 U32 ( .x(n683), .a(Imm[19]) );
	nand2_2 U320 ( .x(n3763), .a(n3482), .b(___cell__39620_net144331) );
	nand2i_4 U3201 ( .x(n2876), .a(n1658), .b(n2802) );
	inv_5 U3203 ( .x(n2944), .a(n3897) );
	nand4_3 U3204 ( .x(n3902), .a(n3901), .b(n3900), .c(n3899), .d(n3898) );
	nand2i_4 U3205 ( .x(n2973), .a(n1626), .b(n2938) );
	nand2i_4 U3207 ( .x(n3944), .a(n1623), .b(n3560) );
	oai211_3 U3208 ( .x(n3110), .a(n630), .b(n718), .c(n3965), .d(n3068) );
	nand2i_2 U321 ( .x(n3438), .a(n1562), .b(n3613) );
	nand2i_4 U3210 ( .x(n3514), .a(n891), .b(n3547) );
	nand4i_4 U3211 ( .x(n3168), .a(n1390), .b(n3974), .c(n3976), .d(n3975) );
	nand2i_4 U3212 ( .x(n3977), .a(n1632), .b(n2994) );
	nand2_5 U3214 ( .x(n3288), .a(n3984), .b(n3175) );
	inv_5 U3215 ( .x(n3204), .a(n3288) );
	nand2_5 U3216 ( .x(n3214), .a(n3985), .b(n3195) );
	nand2i_4 U3217 ( .x(n3210), .a(n1574), .b(n3289) );
	nand4_1 U3218 ( .x(n3990), .a(n3232), .b(n3228), .c(n3225), .d(n3222) );
	nand2i_4 U3219 ( .x(n3991), .a(n1943), .b(___cell__39620_net144303) );
	inv_5 U322 ( .x(n2268), .a(n1730) );
	nand4_1 U3220 ( .x(n1950), .a(n3275), .b(n3271), .c(n3263), .d(n3260) );
	nand3i_3 U3221 ( .x(n3993), .a(n3257), .b(n3256), .c(n3994) );
	nand4_3 U3222 ( .x(n3995), .a(n3287), .b(n3290), .c(n3993), .d(n3282) );
	nand3i_3 U3223 ( .x(n1941), .a(___cell__39620_net144166), .b(n1533), .c(___cell__39620_net143655) );
	inv_5 U3224 ( .x(n2104), .a(n3677) );
	mux2i_3 U3225 ( .x(n2661), .d0(n3383), .sl(n816), .d1(n3386) );
	mux2i_3 U3226 ( .x(n2707), .d0(n3380), .sl(n816), .d1(n3385) );
	mux2i_3 U3227 ( .x(n2797), .d0(n3529), .sl(net149122), .d1(n3534) );
	mux2i_3 U3228 ( .x(n2872), .d0(n3522), .sl(net149122), .d1(n3536) );
	mux2i_3 U3229 ( .x(n3170), .d0(n3515), .sl(net149122), .d1(n3518) );
	nand2_2 U323 ( .x(n1741), .a(n2268), .b(n887) );
	nand2i_4 U3230 ( .x(n1946), .a(IR_opcode_field[0]), .b(N3014) );
	ao221_5 U3232 ( .x(n4070), .a(N361), .b(n977), .c(___cell__39620_net147732),
		.d(n978), .e(n979) );
	nand2_8 U3233 ( .x(n947), .a(___cell__39620_net144312), .b(___cell__39620_net143655) );
	inv_8 U3234 ( .x(n944), .a(n947) );
	inv_10 U3235 ( .x(n3997), .a(n947) );
	nand2i_5 U3236 ( .x(n1455), .a(___cell__39620_net144175), .b(n3995) );
	nor2i_5 U3237 ( .x(n1439), .a(n1440), .b(n1441) );
	nand2i_5 U3238 ( .x(n950), .a(___cell__39620_net143287), .b(n3988) );
	nor3i_5 U3239 ( .x(n967), .a(n3107), .b(n3108), .c(n3105) );
	nand2i_2 U324 ( .x(n2353), .a(n1474), .b(n2139) );
	nor3i_5 U3240 ( .x(n970), .a(n3047), .b(n3048), .c(n3045) );
	and4i_5 U3241 ( .x(n1028), .a(n1345), .b(n1342), .c(n1343), .d(n1344) );
	nor3i_5 U3242 ( .x(n1029), .a(n3006), .b(n3005), .c(n3007) );
	nor3i_5 U3243 ( .x(n951), .a(n1275), .b(n1276), .c(n1277) );
	inv_16 U3244 ( .x(n977), .a(n1596) );
	and4i_5 U3245 ( .x(n980), .a(n2654), .b(n2653), .c(n2657), .d(n2659) );
	nor3i_5 U3246 ( .x(n958), .a(n2096), .b(n2094), .c(n2097) );
	and4i_5 U3247 ( .x(n960), .a(n1059), .b(n1056), .c(n1057), .d(n1058) );
	inv_16 U3248 ( .x(n3057), .a(n1087) );
	aoi21_4 U3249 ( .x(n3161), .a(n1221), .b(n3078), .c(n3158) );
	inv_2 U325 ( .x(n3270), .a(n1474) );
	inv_16 U3250 ( .x(n2837), .a(n1592) );
	nor3i_5 U3251 ( .x(n2881), .a(n2879), .b(n1304), .c(n2880) );
	oai221_5 U3252 ( .x(n2669), .a(n2670), .b(n703), .c(n1234), .d(n4001),
		.e(n2671) );
	oai22_4 U3253 ( .x(n2666), .a(n2667), .b(n784), .c(n2668), .d(___cell__39620_net144406) );
	nand4_2 U3254 ( .x(n2508), .a(n2504), .b(n2509), .c(n2510), .d(n2511) );
	nor3i_5 U3255 ( .x(n1199), .a(n2465), .b(n2463), .c(n2466) );
	aoi21_4 U3256 ( .x(n1200), .a(n662), .b(n2384), .c(n1195) );
	nand2i_5 U3257 ( .x(n2362), .a(n1566), .b(n3752) );
	nand2i_5 U3258 ( .x(n3696), .a(n1694), .b(n3624) );
	oai22_6 U3259 ( .x(___cell__39620_net145444), .a(n784), .b(n696), .c(___cell__39620_net144406),
		.d(n1093) );
	nor2i_1 U326 ( .x(n1179), .a(n534), .b(n4002) );
	inv_16 U3260 ( .x(n1267), .a(n1641) );
	inv_7 U3261 ( .x(n2360), .a(n2238) );
	nand2_8 U3262 ( .x(n1186), .a(n1581), .b(n1576) );
	inv_16 U3263 ( .x(n2024), .a(n670) );
	oai21_6 U3264 ( .x(n2826), .a(n816), .b(n1450), .c(n2808) );
	inv_10 U3265 ( .x(n3662), .a(n1184) );
	inv_10 U3266 ( .x(n3999), .a(n1184) );
	inv_16 U3267 ( .x(n3624), .a(n1169) );
	inv_16 U3268 ( .x(n1064), .a(n1143) );
	aoi222_4 U3269 ( .x(n3169), .a(n3170), .b(n1204), .c(n3171), .d(___cell__39620_net143722),
		.e(n3172), .f(___cell__39620_net143864) );
	inv_4 U327 ( .x(n2206), .a(n3705) );
	inv_16 U3270 ( .x(n1221), .a(n1186) );
	oai221_5 U3271 ( .x(n3078), .a(n3614), .b(n4003), .c(n3611), .d(n1559),
		.e(n3058) );
	nand2i_8 U3272 ( .x(n1588), .a(___cell__39620_net144175), .b(n1589) );
	oai221_5 U3273 ( .x(n2014), .a(n3623), .b(n4004), .c(n3620), .d(n1559),
		.e(n1970) );
	nand2_8 U3274 ( .x(n1574), .a(n1575), .b(n1576) );
	nand2i_5 U3276 ( .x(n3121), .a(n1912), .b(n944) );
	oai221_5 U3277 ( .x(n3041), .a(n3433), .b(n1070), .c(n3600), .d(n1559),
		.e(n3021) );
	nand2i_5 U3278 ( .x(n3099), .a(n1387), .b(n3100) );
	nand2i_5 U3279 ( .x(n3106), .a(n1588), .b(n3041) );
	nor2i_0 U328 ( .x(n2343), .a(n534), .b(n1654) );
	nand2i_5 U3280 ( .x(n1592), .a(___cell__39620_net144175), .b(n1593) );
	inv_16 U3281 ( .x(n1318), .a(n1055) );
	nand3i_5 U3282 ( .x(n3071), .a(n1369), .b(n3072), .c(n3073) );
	aoi22_4 U3283 ( .x(n3080), .a(n1221), .b(n3001), .c(n1191), .d(n3000) );
	nand2i_5 U3284 ( .x(n3037), .a(n1356), .b(n3038) );
	aoi22_4 U3285 ( .x(n3044), .a(n650), .b(n3000), .c(n1221), .d(n3004) );
	nand2i_5 U3286 ( .x(n2984), .a(n1879), .b(n3997) );
	and4i_5 U3287 ( .x(n2950), .a(n2949), .b(n2951), .c(n2948), .d(n2952) );
	nand2i_5 U3288 ( .x(n2964), .a(n1566), .b(n3001) );
	nand2i_6 U3289 ( .x(n2969), .a(n1868), .b(n977) );
	nor2i_1 U329 ( .x(n1163), .a(N1734), .b(___cell__39620_net143710) );
	inv_16 U3290 ( .x(n1197), .a(n1616) );
	nand4i_5 U3291 ( .x(n2846), .a(n1288), .b(n3868), .c(n3870), .d(n3869) );
	inv_16 U3292 ( .x(n4000), .a(n946) );
	nand2i_5 U3293 ( .x(n2885), .a(n1855), .b(n1987) );
	nand2i_5 U3294 ( .x(n2886), .a(n1854), .b(n3662) );
	nand3i_5 U3295 ( .x(n2893), .a(n1310), .b(n2894), .c(n2895) );
	oai211_5 U3296 ( .x(n2849), .a(n3629), .b(n1043), .c(n2765), .d(n3859) );
	nand2_8 U3297 ( .x(n1626), .a(n1436), .b(___cell__39620_net147732) );
	nand2i_6 U3298 ( .x(n2832), .a(n1574), .b(n3752) );
	nand2i_5 U3299 ( .x(n2833), .a(n1566), .b(n3289) );
	inv_2 U330 ( .x(n4002), .a(n766) );
	inv_16 U3300 ( .x(___cell__39620_net143722), .a(___cell__39620_net144406) );
	nand2_5 U3301 ( .x(n2757), .a(n513), .b(n502) );
	nand2_5 U3302 ( .x(n2758), .a(n2797), .b(n1267) );
	oai221_5 U3303 ( .x(n2557), .a(n1315), .b(n1043), .c(n3426), .d(n1072),
		.e(n1806) );
	nand2i_5 U3304 ( .x(n2686), .a(n1166), .b(n2733) );
	ao222_5 U3305 ( .x(n2706), .a(n2707), .b(n2024), .c(n745), .d(___cell__39620_net145617),
		.e(n2708), .f(n2022) );
	oai221_5 U3306 ( .x(n2532), .a(n3420), .b(n4003), .c(n1300), .d(n1565),
		.e(n1807) );
	inv_16 U3307 ( .x(n1191), .a(n1588) );
	nand2_5 U3308 ( .x(n2664), .a(n2708), .b(n1267) );
	inv_6 U3309 ( .x(n1234), .a(n3821) );
	nand2_8 U3310 ( .x(n1658), .a(n1429), .b(___cell__39620_net147732) );
	nand2_8 U3311 ( .x(n4001), .a(n1429), .b(___cell__39620_net147732) );
	nand2i_8 U3312 ( .x(___cell__39620_net144406), .a(___cell__39620_net144175),
		.b(n1650) );
	nand2i_5 U3313 ( .x(n2597), .a(n1795), .b(n3662) );
	nor2i_5 U3314 ( .x(n1225), .a(n1085), .b(n1211) );
	nand2i_5 U3315 ( .x(n2575), .a(n1220), .b(n2576) );
	nand2i_4 U3316 ( .x(n2539), .a(n784), .b(n3796) );
	oai22_6 U3317 ( .x(n2490), .a(n1637), .b(n1122), .c(n1626), .d(n1120) );
	aoai211_5 U3318 ( .x(n2528), .a(n1267), .b(n2570), .c(n3809), .d(___cell__39620_net144345) );
	nand2i_5 U3319 ( .x(n2516), .a(n1779), .b(___cell__39620_net145508) );
	oai22_1 U332 ( .x(n2838), .a(n679), .b(n4026), .c(n1602), .d(n4002) );
	nand2i_5 U3320 ( .x(n2465), .a(n1767), .b(n3997) );
	nor2i_5 U3321 ( .x(n1203), .a(n1204), .b(n1205) );
	nand2i_5 U3322 ( .x(n2445), .a(n703), .b(n2391) );
	aoi22_4 U3323 ( .x(n2422), .a(n1318), .b(n2384), .c(n1095), .d(n2423) );
	aoi21_6 U3325 ( .x(n2368), .a(n2024), .b(n2371), .c(n1180) );
	nand2i_6 U3326 ( .x(n2370), .a(n1626), .b(n3711) );
	inv_6 U3327 ( .x(n2359), .a(n2192) );
	nand2i_6 U3328 ( .x(n2332), .a(n1658), .b(___cell__39620_net147278) );
	nand3i_5 U3329 ( .x(n1077), .a(n1614), .b(n810), .c(___cell__39620_net144355) );
	exnor2_1 U333 ( .x(n1496), .a(n815), .b(n692) );
	aoi21_4 U3330 ( .x(n2246), .a(n2022), .b(n2247), .c(n2248) );
	nand2i_5 U3331 ( .x(n2171), .a(n1124), .b(n2172) );
	aoi22_4 U3332 ( .x(n2164), .a(n2161), .b(___cell__39620_net147791), .c(n1095),
		.d(n2165) );
	inv_16 U3333 ( .x(___cell__39620_net143864), .a(n784) );
	inv_16 U3334 ( .x(n1204), .a(n4001) );
	oai21_5 U3335 ( .x(n2103), .a(n703), .b(n2104), .c(n2105) );
	nand2i_4 U3336 ( .x(n2101), .a(n1626), .b(n2059) );
	aoi21_5 U3337 ( .x(n2098), .a(n502), .b(n2099), .c(n1106) );
	nand2i_4 U3338 ( .x(n2034), .a(n784), .b(n2064) );
	nor2i_1 U334 ( .x(n1284), .a(n1285), .b(n690) );
	aoi21_5 U3340 ( .x(n3195), .a(n1256), .b(n3196), .c(n3197) );
	nand2_8 U3341 ( .x(n1641), .a(n1428), .b(___cell__39620_net143326) );
	inv_16 U3342 ( .x(___cell__39620_net144345), .a(net149122) );
	inv_16 U3343 ( .x(n1657), .a(n917) );
	oai211_5 U3344 ( .x(n2238), .a(n3430), .b(n815), .c(n3431), .d(n3432) );
	inv_16 U3345 ( .x(n2139), .a(n1536) );
	inv_12 U3346 ( .x(___cell__39620_net147791), .a(___cell__39620_net143658) );
	and2_8 U3347 ( .x(n1422), .a(n1197), .b(n1423) );
	nand4i_5 U3348 ( .x(n1988), .a(n1041), .b(n3634), .c(n3633), .d(n3632) );
	inv_16 U3349 ( .x(n1095), .a(n1166) );
	inv_2 U335 ( .x(n1285), .a(n1495) );
	nand4i_5 U3350 ( .x(n1992), .a(n1048), .b(n3661), .c(n3660), .d(n3659) );
	inv_16 U3351 ( .x(n1987), .a(n1077) );
	nand2i_8 U3352 ( .x(n1143), .a(___cell__39620_net144175), .b(n1710) );
	nand2i_8 U3353 ( .x(___cell__39620_net143693), .a(n1618), .b(___cell__39620_net143326) );
	oai211_4 U3354 ( .x(n2023), .a(n3452), .b(n1625), .c(n3590), .d(n1994) );
	inv_16 U3355 ( .x(n1085), .a(n703) );
	nand2i_5 U3356 ( .x(n4003), .a(reg_out_B[3]), .b(n815) );
	nand2i_4 U3357 ( .x(n4004), .a(reg_out_B[3]), .b(n815) );
	nand2i_8 U3358 ( .x(n1559), .a(n815), .b(reg_out_B[3]) );
	aoi22_4 U3359 ( .x(n3058), .a(n1971), .b(n3059), .c(n1330), .d(n1965) );
	exnor2_1 U336 ( .x(n1495), .a(n891), .b(n692) );
	aoi22_4 U3360 ( .x(n1970), .a(n1971), .b(n1972), .c(n1330), .d(n1069) );
	oai221_4 U3361 ( .x(n2054), .a(n3433), .b(n1559), .c(n3600), .d(n1562),
		.e(n1967) );
	nand2i_8 U3362 ( .x(n1055), .a(___cell__39620_net144345), .b(___cell__39620_net144347) );
	nand4i_5 U3363 ( .x(n1380), .a(n1348), .b(n3960), .c(n3959), .d(n3958) );
	oai221_4 U3365 ( .x(n3112), .a(n3355), .b(n1635), .c(n849), .d(n727), .e(n3070) );
	nand2i_5 U3366 ( .x(n3100), .a(n702), .b(n3076) );
	oai211_5 U3367 ( .x(n3075), .a(n3515), .b(___cell__39620_net144345), .c(n3972),
		.d(n3971) );
	oai221_5 U3368 ( .x(n3000), .a(n3439), .b(n4003), .c(n747), .d(n1559),
		.e(n2980) );
	nor2i_5 U3369 ( .x(n1332), .a(n1333), .b(n1334) );
	nand2i_2 U337 ( .x(n3757), .a(n2339), .b(n3756) );
	nand2i_5 U3370 ( .x(n3953), .a(n4007), .b(n3646) );
	oai211_4 U3371 ( .x(n3051), .a(n3452), .b(n4008), .c(n3957), .d(n3032) );
	nand2i_5 U3372 ( .x(n3072), .a(n702), .b(n3963) );
	nand2i_6 U3373 ( .x(n3073), .a(n4001), .b(n3040) );
	oai211_4 U3374 ( .x(n3076), .a(n3413), .b(n1451), .c(n3970), .d(n3969) );
	nand4i_5 U3375 ( .x(n3001), .a(n1321), .b(n3934), .c(n3933), .d(n3932) );
	nand2i_5 U3376 ( .x(n3936), .a(n1072), .b(n3628) );
	nand2i_6 U3377 ( .x(n3935), .a(n1607), .b(n3774) );
	nand4i_5 U3378 ( .x(n1339), .a(n1314), .b(n3909), .c(n3908), .d(n3907) );
	oai221_4 U3379 ( .x(n3054), .a(n3366), .b(n1632), .c(n511), .d(n1636),
		.e(n3035) );
	nand2_2 U338 ( .x(n2339), .a(n2340), .b(n2341) );
	nand2i_5 U3380 ( .x(n3038), .a(___cell__39620_net144406), .b(n3963) );
	oai211_5 U3381 ( .x(n3040), .a(n499), .b(___cell__39620_net144345), .c(n3961),
		.d(n3962) );
	nand4i_5 U3382 ( .x(n3004), .a(n1312), .b(n3906), .c(n3905), .d(n3904) );
	nand4i_5 U3383 ( .x(n1308), .a(n1301), .b(n3884), .c(n3883), .d(n3882) );
	ao22_6 U3385 ( .x(n2949), .a(n662), .b(n2846), .c(n1318), .d(n1308) );
	nand4i_5 U3386 ( .x(n2859), .a(n1286), .b(n3867), .c(n3866), .d(n3865) );
	aoi21_5 U3387 ( .x(n2917), .a(n662), .b(n2849), .c(n1316) );
	nor2i_5 U3388 ( .x(n1317), .a(n1318), .b(n1319) );
	nand2_8 U3389 ( .x(___cell__39620_net143653), .a(IR_opcode_field[1]), .b(IR_opcode_field[0]) );
	inv_4 U339 ( .x(n3341), .a(n3470) );
	nand2i_6 U3390 ( .x(n1616), .a(net149122), .b(___cell__39620_net143785) );
	nor2i_5 U3391 ( .x(n1288), .a(n1289), .b(n1290) );
	nand2i_5 U3392 ( .x(n3868), .a(n4006), .b(n3648) );
	nand2i_6 U3393 ( .x(n3870), .a(n4005), .b(n3646) );
	nand2i_8 U3394 ( .x(n1182), .a(___cell__39620_net144345), .b(___cell__39620_net143785) );
	nand2i_6 U3395 ( .x(n1166), .a(net149120), .b(___cell__39620_net144347) );
	oai211_5 U3396 ( .x(n2863), .a(n3611), .b(n1565), .c(n3850), .d(n2718) );
	nand2i_6 U3397 ( .x(n2892), .a(n3889), .b(n1217) );
	oai211_5 U3399 ( .x(n2911), .a(n3460), .b(n4008), .c(n3876), .d(n2889) );
	inv_2 U34 ( .x(n596), .a(n886) );
	oai211_1 U340 ( .x(n2337), .a(n3341), .b(___cell__39620_net144317), .c(n3342),
		.d(n2163) );
	or2_8 U3400 ( .x(n4005), .a(n891), .b(net149167) );
	inv_16 U3401 ( .x(n2193), .a(n1116) );
	nand2i_6 U3402 ( .x(n2856), .a(n3875), .b(n1217) );
	oai211_5 U3403 ( .x(n2192), .a(n3436), .b(n815), .c(n3437), .d(n3438) );
	nand2i_6 U3404 ( .x(n3864), .a(net149120), .b(n1431) );
	nand2i_5 U3406 ( .x(n2769), .a(n1055), .b(n2733) );
	aoi21_5 U3407 ( .x(n2780), .a(n1714), .b(n2781), .c(n1258) );
	aoi21_4 U3408 ( .x(n2778), .a(n504), .b(n2779), .c(n1255) );
	inv_10 U3409 ( .x(n2746), .a(n2863) );
	nor2i_1 U341 ( .x(n1270), .a(N1700), .b(___cell__39620_net143660) );
	inv_10 U3410 ( .x(n1298), .a(n2902) );
	oai22_6 U3411 ( .x(n2723), .a(___cell__39620_net143710), .b(n1820), .c(___cell__39620_net143658),
		.d(n2720) );
	nand2_5 U3412 ( .x(n2756), .a(n2710), .b(n2022) );
	nand2i_4 U3413 ( .x(n4006), .a(net149167), .b(n891) );
	nand2i_4 U3414 ( .x(n4007), .a(net149167), .b(n891) );
	nand2i_8 U3415 ( .x(n1806), .a(n4140), .b(net149167) );
	nand4_3 U3417 ( .x(n3835), .a(n3834), .b(n3833), .c(n3832), .d(n3831) );
	nor2i_8 U3418 ( .x(n1237), .a(N1853), .b(n946) );
	nand2_8 U3419 ( .x(n1807), .a(n1728), .b(reg_out_B[3]) );
	inv_2 U342 ( .x(n1272), .a(N1865) );
	inv_7 U3420 ( .x(n1429), .a(n1653) );
	nand2i_5 U3421 ( .x(n2601), .a(n1182), .b(n2473) );
	nand2i_5 U3422 ( .x(n2576), .a(n1588), .b(n3422) );
	oai21_5 U3423 ( .x(n2582), .a(n621), .b(n2583), .c(n2584) );
	oai211_5 U3424 ( .x(n2473), .a(n3427), .b(n1602), .c(n3428), .d(n3429) );
	oai21_6 U3425 ( .x(n2423), .a(n3421), .b(n4005), .c(n3572) );
	nand2_8 U3426 ( .x(n3571), .a(n1728), .b(n1565) );
	nand2i_8 U3427 ( .x(n1122), .a(n1635), .b(n883) );
	nand2i_8 U3428 ( .x(n1120), .a(n718), .b(n4130) );
	aoi21_6 U3429 ( .x(n2503), .a(N1757), .b(___cell__39620_net145150), .c(n1207) );
	nor2_1 U343 ( .x(n1271), .a(n947), .b(n1272) );
	nand2i_6 U3430 ( .x(n2513), .a(n1778), .b(n1987) );
	nor2i_8 U3431 ( .x(n1196), .a(n1197), .b(n1198) );
	nand2i_5 U3433 ( .x(n2446), .a(n1566), .b(n2492) );
	nor2i_8 U3434 ( .x(n1189), .a(N1858), .b(n946) );
	oai21_6 U3436 ( .x(n2319), .a(n694), .b(n3735), .c(n2301) );
	oai211_4 U3437 ( .x(n2168), .a(n891), .b(n3506), .c(n3507), .d(n3508) );
	inv_16 U3438 ( .x(n1646), .a(n692) );
	or2_8 U3439 ( .x(n4008), .a(n637), .b(net149120) );
	nor2i_1 U344 ( .x(n2811), .a(n891), .b(n1646) );
	nand2i_5 U3440 ( .x(n2256), .a(n670), .b(n3702) );
	oai211_5 U3441 ( .x(n2089), .a(n3439), .b(n1562), .c(n3440), .d(n3441) );
	nand2i_5 U3442 ( .x(n2172), .a(n1182), .b(n2043) );
	nand2i_6 U3443 ( .x(n2190), .a(n3709), .b(n1217) );
	nand4i_5 U3444 ( .x(n2090), .a(n1068), .b(n3672), .c(n3671), .d(n3670) );
	nand4i_5 U3445 ( .x(n1993), .a(n1044), .b(n3643), .c(n3642), .d(n3641) );
	nand4i_5 U3446 ( .x(n2043), .a(n1071), .b(n3675), .c(n3674), .d(n3673) );
	nand2i_5 U3447 ( .x(n2145), .a(n1588), .b(n2090) );
	nor2i_8 U3448 ( .x(n1096), .a(N1738), .b(___cell__39620_net143710) );
	nor2i_8 U3449 ( .x(n1099), .a(N1837), .b(n946) );
	inv_2 U345 ( .x(n1274), .a(N1799) );
	oai221_4 U3450 ( .x(n2093), .a(n3614), .b(n1559), .c(n3611), .d(n1562),
		.e(n1963) );
	nand2_8 U3451 ( .x(n2060), .a(n3677), .b(___cell__39620_net143722) );
	nand2i_6 U3452 ( .x(n2061), .a(n1626), .b(n3583) );
	oai21_5 U3453 ( .x(n2062), .a(n784), .b(n870), .c(n2063) );
	nand2i_6 U3454 ( .x(n2009), .a(n1457), .b(n2139) );
	aoi21_5 U3455 ( .x(n3175), .a(n1256), .b(n3176), .c(n3177) );
	nand2i_8 U3456 ( .x(n1040), .a(n759), .b(n1553) );
	nand2i_6 U3457 ( .x(n1446), .a(n1535), .b(n1528) );
	aoi21_6 U3458 ( .x(n1430), .a(n694), .b(n1431), .c(n1432) );
	nand2i_6 U3459 ( .x(n1639), .a(n1640), .b(n676) );
	nor2_1 U346 ( .x(n1273), .a(n1077), .b(n1274) );
	oai211_5 U3460 ( .x(n3196), .a(n3345), .b(n1546), .c(n3349), .d(n3350) );
	inv_16 U3461 ( .x(n1643), .a(n4011) );
	inv_16 U3462 ( .x(n1066), .a(n4010) );
	inv_16 U3463 ( .x(n1714), .a(n1635) );
	nand2i_6 U3465 ( .x(n3538), .a(n501), .b(n3627) );
	nor2i_6 U3466 ( .x(n1041), .a(n1042), .b(n1043) );
	nand2i_5 U3467 ( .x(n3634), .a(n1608), .b(n3628) );
	nand2i_5 U3468 ( .x(n3633), .a(n4007), .b(n3538) );
	nand2i_6 U3469 ( .x(n3632), .a(n1607), .b(n2766) );
	nand3_4 U347 ( .x(n1165), .a(n3754), .b(n665), .c(n2344) );
	nor2i_6 U3470 ( .x(n1360), .a(n1361), .b(n4005) );
	nand2i_5 U3471 ( .x(n3967), .a(n4007), .b(n3537) );
	nand2i_6 U3472 ( .x(n3966), .a(n1607), .b(n2722) );
	nand2i_5 U3473 ( .x(n3651), .a(n1608), .b(n3646) );
	nand2i_6 U3474 ( .x(n3649), .a(n1607), .b(n3648) );
	nor2i_5 U3475 ( .x(n1390), .a(n1391), .b(n1392) );
	nand2i_5 U3476 ( .x(n3974), .a(n4010), .b(n4142) );
	nand2i_6 U3477 ( .x(n3976), .a(n4008), .b(n2181) );
	nand2i_6 U3478 ( .x(n1625), .a(n694), .b(n891) );
	inv_6 U3479 ( .x(n3515), .a(n3512) );
	nand2i_2 U348 ( .x(n2137), .a(n1064), .b(n3698) );
	nand2i_6 U3480 ( .x(n3622), .a(n3621), .b(n3598) );
	nand2i_6 U3481 ( .x(n1972), .a(n3585), .b(n3617) );
	nor2i_6 U3482 ( .x(n1348), .a(n1349), .b(n1043) );
	nand2i_5 U3483 ( .x(n3960), .a(n1608), .b(n3655) );
	nand2i_5 U3484 ( .x(n3959), .a(n4007), .b(n3658) );
	nand2i_6 U3485 ( .x(n3958), .a(n1607), .b(n2677) );
	nand2i_5 U3486 ( .x(n1701), .a(___cell__39620_net144175), .b(n1939) );
	nand2i_6 U3487 ( .x(n3022), .a(n3585), .b(n3801) );
	aoi22_4 U3488 ( .x(n3068), .a(n1066), .b(n2991), .c(n1391), .d(n3069) );
	nand2i_6 U3489 ( .x(n3972), .a(n4008), .b(n2927) );
	nor2i_1 U349 ( .x(n2108), .a(n1451), .b(___cell__39620_net144406) );
	nand2i_5 U3490 ( .x(n3971), .a(n4010), .b(n3560) );
	aoi21_5 U3491 ( .x(n2980), .a(n1971), .b(n2981), .c(n1329) );
	nand2i_6 U3492 ( .x(n1608), .a(n891), .b(net149167) );
	nand2i_6 U3493 ( .x(n3790), .a(n751), .b(n3789) );
	nor2i_5 U3494 ( .x(n1321), .a(n1177), .b(n1322) );
	nand2i_5 U3495 ( .x(n3934), .a(n1070), .b(n3619) );
	nand2i_6 U3496 ( .x(n3932), .a(n1562), .b(n2763) );
	inv_16 U3497 ( .x(n1147), .a(n1608) );
	nand2i_6 U3498 ( .x(n3774), .a(n751), .b(n3773) );
	nor2i_8 U3499 ( .x(n1314), .a(n1147), .b(n1315) );
	inv_5 U35 ( .x(n640), .a(n638) );
	nor2_1 U350 ( .x(n2109), .a(n784), .b(n694) );
	nand2i_6 U3500 ( .x(n3909), .a(n4005), .b(n3537) );
	nand2i_5 U3501 ( .x(n3908), .a(n4006), .b(n3638) );
	nand2i_6 U3502 ( .x(n3907), .a(n1607), .b(n3764) );
	nand2i_6 U3503 ( .x(n3962), .a(n4008), .b(n2783) );
	nor2i_5 U3504 ( .x(n1312), .a(n1177), .b(n1313) );
	nor2i_5 U3505 ( .x(n1301), .a(n1147), .b(n1302) );
	nand2i_5 U3506 ( .x(n3883), .a(n1072), .b(n3655) );
	nand2i_6 U3507 ( .x(n3882), .a(n1607), .b(n3744) );
	nor2i_5 U3508 ( .x(n1299), .a(n1177), .b(n1300) );
	nand2i_6 U3509 ( .x(n3880), .a(n1565), .b(n3602) );
	aoi222_1 U351 ( .x(n2134), .a(n2109), .b(n2135), .c(n2108), .d(n2136),
		.e(reg_out_B[6]), .f(n2137) );
	nand2i_6 U3510 ( .x(n3879), .a(n1562), .b(n2673) );
	nand2i_6 U3511 ( .x(n2998), .a(n1505), .b(n2139) );
	nor2i_5 U3512 ( .x(n1286), .a(n1177), .b(n1287) );
	nand2i_5 U3513 ( .x(n3867), .a(n1070), .b(n685) );
	nand2i_6 U3514 ( .x(n2960), .a(n1503), .b(n2139) );
	oai211_4 U3515 ( .x(n3897), .a(n3553), .b(n4008), .c(n3896), .d(n2926) );
	nand2i_5 U3516 ( .x(n2972), .a(n670), .b(n3902) );
	nand2i_5 U3517 ( .x(n3877), .a(n1634), .b(n3020) );
	nand2i_6 U3518 ( .x(n2935), .a(n1502), .b(n2139) );
	oai211_5 U3519 ( .x(n3887), .a(n3522), .b(___cell__39620_net144345), .c(n3886),
		.d(n3885) );
	aoi21_1 U352 ( .x(n2138), .a(n2139), .b(n2140), .c(n1114) );
	nand2i_6 U3520 ( .x(n3913), .a(n1417), .b(n530) );
	nand2i_5 U3521 ( .x(n3857), .a(n4004), .b(n1972) );
	nand2i_5 U3522 ( .x(n2915), .a(n1861), .b(___cell__39620_net145150) );
	aoi21_5 U3523 ( .x(n2718), .a(n1177), .b(n2719), .c(n2630) );
	inv_6 U3525 ( .x(n3529), .a(n3526) );
	nand2i_6 U3526 ( .x(n3872), .a(n4008), .b(n3069) );
	aoi22_4 U3527 ( .x(n2889), .a(n1391), .b(n2890), .c(n1066), .d(n2783) );
	nand2i_6 U3528 ( .x(n2766), .a(n751), .b(n3631) );
	nand2_8 U3529 ( .x(n1623), .a(n694), .b(n891) );
	inv_2 U353 ( .x(n2140), .a(n1464) );
	nand2i_5 U3530 ( .x(n3845), .a(n1070), .b(n3022) );
	nand2i_6 U3531 ( .x(n3537), .a(n3565), .b(n3627) );
	nand2i_6 U3532 ( .x(n3756), .a(n816), .b(n3755) );
	nand2i_5 U3533 ( .x(n3437), .a(n1070), .b(n1966) );
	inv_16 U3534 ( .x(___cell__39620_net144517), .a(___cell__39620_net144374) );
	inv_16 U3536 ( .x(n1391), .a(n1623) );
	nand4i_5 U3537 ( .x(n1431), .a(n1282), .b(n3861), .c(n2804), .d(n3863) );
	oai21_5 U3538 ( .x(n3365), .a(n3366), .b(n815), .c(n3367) );
	oai21_6 U3539 ( .x(n2781), .a(n2429), .b(n536), .c(n3400) );
	exnor2_1 U354 ( .x(n1464), .a(reg_out_B[6]), .b(n922) );
	nor2i_5 U3540 ( .x(n1258), .a(n1249), .b(n1259) );
	nor2i_8 U3541 ( .x(n1255), .a(n1256), .b(n1257) );
	aoi22_4 U3542 ( .x(n2782), .a(n1391), .b(n2783), .c(n1066), .d(n2784) );
	aoi21_4 U3544 ( .x(n2721), .a(n2676), .b(n2722), .c(n2634) );
	nand2i_5 U3545 ( .x(n3855), .a(n1608), .b(n3764) );
	nand2i_5 U3546 ( .x(n3846), .a(n1608), .b(n3744) );
	nand2i_6 U3547 ( .x(n2744), .a(n1816), .b(n530) );
	aoi21_4 U3548 ( .x(n2632), .a(n1147), .b(n2633), .c(n2634) );
	nand2i_5 U3549 ( .x(n3838), .a(n4007), .b(n3790) );
	nor2i_1 U355 ( .x(n1114), .a(n1115), .b(n690) );
	nand2_4 U3550 ( .x(n3834), .a(n504), .b(n2373) );
	nand2i_6 U3552 ( .x(n2673), .a(n3585), .b(n3742) );
	nand2i_6 U3553 ( .x(n2763), .a(n3585), .b(n3772) );
	nand2i_6 U3554 ( .x(n2719), .a(n3585), .b(n3762) );
	nand2i_6 U3555 ( .x(n3840), .a(n1797), .b(n530) );
	nand2i_5 U3556 ( .x(n2591), .a(n2588), .b(___cell__39620_net147791) );
	nand2_3 U3557 ( .x(n3814), .a(n1714), .b(n2373) );
	nand2i_8 U3558 ( .x(n1645), .a(n1560), .b(n883) );
	nand2i_6 U3559 ( .x(n3428), .a(n4140), .b(n1147) );
	inv_2 U356 ( .x(n1115), .a(n1463) );
	nand2i_6 U3560 ( .x(n3429), .a(n1043), .b(n3790) );
	nand2i_6 U3561 ( .x(n3804), .a(n1771), .b(n530) );
	nand2i_6 U3562 ( .x(n3744), .a(n751), .b(n3743) );
	oai21_6 U3563 ( .x(n3778), .a(n1587), .b(n1642), .c(n3777) );
	nand2i_6 U3564 ( .x(n2410), .a(n2411), .b(n1217) );
	inv_10 U3565 ( .x(n1555), .a(n1554) );
	inv_6 U3566 ( .x(n3731), .a(n3730) );
	nand2i_6 U3567 ( .x(n2397), .a(n1476), .b(n2139) );
	nand2i_6 U3568 ( .x(n3508), .a(n1607), .b(n3658) );
	oai22_6 U3569 ( .x(n2148), .a(n784), .b(n1120), .c(___cell__39620_net144406),
		.d(n1122) );
	nand2i_2 U357 ( .x(n2144), .a(n1574), .b(n2089) );
	inv_16 U3570 ( .x(n1177), .a(n1559) );
	inv_16 U3571 ( .x(n1683), .a(n4008) );
	nand2i_6 U3572 ( .x(n2322), .a(n1472), .b(n2139) );
	nand2i_6 U3573 ( .x(n2292), .a(n1470), .b(n2139) );
	nand2i_6 U3574 ( .x(n3441), .a(n815), .b(n3683) );
	inv_16 U3575 ( .x(n1656), .a(n912) );
	nand2i_6 U3576 ( .x(n3672), .a(n1562), .b(n3619) );
	nor2i_8 U3577 ( .x(n1044), .a(n1045), .b(n4005) );
	nand2i_5 U3578 ( .x(n3643), .a(n1608), .b(n3537) );
	nand2i_5 U3579 ( .x(n3642), .a(n1072), .b(n1361) );
	nand3_2 U358 ( .x(n2099), .a(n2081), .b(n3685), .c(n2084) );
	nand2i_6 U3580 ( .x(n3641), .a(n1607), .b(n3638) );
	nand2i_6 U3581 ( .x(n3674), .a(n1607), .b(n3628) );
	oai22_6 U3582 ( .x(n2136), .a(n1642), .b(n1656), .c(n915), .d(n1657) );
	nor2i_5 U3583 ( .x(n1065), .a(n1066), .b(n1067) );
	nand2i_5 U3584 ( .x(n3680), .a(n4010), .b(n2181) );
	nand2i_6 U3585 ( .x(n2048), .a(n1459), .b(n2139) );
	inv_16 U3586 ( .x(n1529), .a(n904) );
	nand2i_6 U3587 ( .x(n3580), .a(n1623), .b(n4142) );
	inv_7 U3588 ( .x(n1553), .a(n1157) );
	oai21_6 U3589 ( .x(n1836), .a(n1642), .b(n1646), .c(n1837) );
	nand2i_2 U359 ( .x(n2150), .a(n670), .b(n2099) );
	inv_16 U3590 ( .x(n3591), .a(n1642) );
	nand2i_5 U3591 ( .x(n1432), .a(n3233), .b(n3234) );
	nand3i_5 U3592 ( .x(n3182), .a(n1416), .b(n3183), .c(n3184) );
	nor2i_5 U3593 ( .x(n1176), .a(n1177), .b(n1178) );
	aoi21_5 U3594 ( .x(n2338), .a(n1971), .b(n2184), .c(n1174) );
	nand2i_6 U3595 ( .x(n3416), .a(n1655), .b(n3592) );
	nand2_8 U3596 ( .x(n3349), .a(n1691), .b(n628) );
	nand2i_6 U3597 ( .x(n3350), .a(n1656), .b(n883) );
	nand2_8 U3598 ( .x(n1690), .a(n1691), .b(n504) );
	buf_16 U3599 ( .x(n4011), .a(n1631) );
	inv_8 U36 ( .x(net156363), .a(___cell__39620_net143997) );
	nor2_1 U360 ( .x(n1117), .a(n4002), .b(___cell__39620_net143735) );
	aoi22_4 U3600 ( .x(n2334), .a(n1289), .b(n2080), .c(n2335), .d(n636) );
	nand2_8 U3601 ( .x(n3342), .a(n1686), .b(n628) );
	nand2i_6 U3603 ( .x(n3412), .a(n1644), .b(n3592) );
	nand2i_8 U3604 ( .x(n3638), .a(n3389), .b(n3627) );
	nand2i_8 U3605 ( .x(n3655), .a(n3486), .b(n3627) );
	nand2_3 U3606 ( .x(n3980), .a(n504), .b(n2187) );
	nand2_3 U3607 ( .x(n3979), .a(n1714), .b(n2000) );
	oai22_6 U3608 ( .x(n3356), .a(n915), .b(n1656), .c(n3357), .d(n815) );
	oai22_6 U3609 ( .x(n3530), .a(n891), .b(n3294), .c(n1651), .d(n1656) );
	inv_2 U361 ( .x(n3505), .a(n2045) );
	nand2_8 U3610 ( .x(n3817), .a(n3311), .b(n855) );
	nand2_8 U3611 ( .x(n3617), .a(n3556), .b(n855) );
	inv_16 U3612 ( .x(n1586), .a(n901) );
	nand2i_6 U3613 ( .x(n2677), .a(n751), .b(n3802) );
	oai22_6 U3614 ( .x(n3036), .a(n1573), .b(n1629), .c(n1569), .d(n825) );
	nand2_8 U3615 ( .x(n2991), .a(n3567), .b(n3568) );
	nand2_8 U3616 ( .x(n3069), .a(n3361), .b(n3362) );
	nand2_8 U3617 ( .x(n2927), .a(n3297), .b(n3298) );
	nor2i_5 U3618 ( .x(n1329), .a(n1330), .b(n1331) );
	inv_10 U3619 ( .x(n1605), .a(n3576) );
	mux2i_1 U362 ( .x(n2157), .d0(n3546), .sl(n816), .d1(n3442) );
	nand2_6 U3620 ( .x(n3033), .a(n3363), .b(n3364) );
	oai22_6 U3621 ( .x(n2852), .a(n1629), .b(n1649), .c(n1579), .d(n881) );
	nand2_8 U3622 ( .x(n2854), .a(n3372), .b(n3373) );
	inv_16 U3623 ( .x(n1571), .a(n644) );
	nand2_8 U3624 ( .x(n2783), .a(n3300), .b(n3301) );
	oai22_6 U3625 ( .x(n2851), .a(n1571), .b(n881), .c(n1629), .d(n1644) );
	inv_7 U3626 ( .x(n1287), .a(n2981) );
	nand2i_5 U3627 ( .x(n2629), .a(n1156), .b(n1558) );
	aoi22_6 U3628 ( .x(n2926), .a(n1066), .b(n2927), .c(___cell__39620_net144517),
		.d(n2854) );
	nand2i_5 U3629 ( .x(n3901), .a(n1635), .b(n2995) );
	nor2_1 U363 ( .x(n1118), .a(n1087), .b(n4042) );
	oai22_6 U3630 ( .x(n3020), .a(n1629), .b(n1656), .c(n1563), .d(n881) );
	nand2i_6 U3631 ( .x(n2633), .a(n1605), .b(n3725) );
	nand2i_6 U3632 ( .x(n3888), .a(n1851), .b(n530) );
	nand2_8 U3633 ( .x(n2784), .a(n3376), .b(n3377) );
	nand2_6 U3634 ( .x(n2890), .a(n3295), .b(n3296) );
	nand2i_6 U3635 ( .x(n3569), .a(n4140), .b(n1289) );
	oai22_6 U3636 ( .x(n3535), .a(n891), .b(n3306), .c(n1573), .d(n1651) );
	buf_16 U3639 ( .x(n4013), .a(n1622) );
	inv_2 U364 ( .x(n1113), .a(N1869) );
	nor2i_5 U3640 ( .x(n1282), .a(n1147), .b(n1283) );
	nand2i_6 U3641 ( .x(n3863), .a(n1644), .b(n811) );
	nand2i_6 U3642 ( .x(n3367), .a(n1578), .b(n3592) );
	nand2i_6 U3643 ( .x(n3400), .a(n1529), .b(n3584) );
	nor2i_5 U3644 ( .x(n1248), .a(n1249), .b(n1250) );
	oai21_6 U3645 ( .x(n2649), .a(n4125), .b(n1148), .c(n3453) );
	nand2_8 U3646 ( .x(n3742), .a(n3351), .b(n855) );
	nand2_8 U3647 ( .x(n3772), .a(n3332), .b(n855) );
	nand2i_6 U3648 ( .x(n2262), .a(n3565), .b(n3566) );
	nand2i_6 U3649 ( .x(n2277), .a(n501), .b(n3501) );
	nor2_1 U365 ( .x(n1112), .a(n947), .b(n1113) );
	nand2i_6 U3650 ( .x(n3791), .a(n1760), .b(n1063) );
	nand2i_6 U3651 ( .x(n3786), .a(n4140), .b(n2458) );
	oai211_5 U3652 ( .x(n2305), .a(n506), .b(n1546), .c(n3401), .d(n3402) );
	nand2i_6 U3653 ( .x(n3718), .a(n1580), .b(n3591) );
	nand2_8 U3654 ( .x(n3407), .a(n1691), .b(n908) );
	nand2i_6 U3655 ( .x(n3408), .a(n1573), .b(n883) );
	nand2i_6 U3656 ( .x(n3721), .a(n1578), .b(n811) );
	aoi21_4 U3657 ( .x(n2276), .a(n1289), .b(n2277), .c(n1146) );
	nand2i_6 U3658 ( .x(n3722), .a(n1580), .b(n3594) );
	nor2i_1 U366 ( .x(n1111), .a(N1737), .b(___cell__39620_net143710) );
	nand2_8 U3660 ( .x(n3398), .a(n1686), .b(n908) );
	nand2i_6 U3661 ( .x(n3399), .a(n1573), .b(n928) );
	aoi21_6 U3662 ( .x(n2065), .a(n2066), .b(n634), .c(n2067) );
	nand2i_6 U3663 ( .x(n3733), .a(n1219), .b(n811) );
	aoi21_4 U3664 ( .x(n2261), .a(n1289), .b(n2262), .c(n1151) );
	nor2i_8 U3665 ( .x(n1109), .a(n686), .b(n1091) );
	inv_16 U3666 ( .x(n1644), .a(n922) );
	nand2i_6 U3667 ( .x(n2080), .a(n1605), .b(n3577) );
	nor2i_8 U3668 ( .x(n1090), .a(n634), .b(n1091) );
	nand2i_8 U3669 ( .x(n1687), .a(n1546), .b(n504) );
	nand2i_2 U367 ( .x(n3103), .a(n1512), .b(n2139) );
	nand2i_6 U3670 ( .x(n3183), .a(n1682), .b(n1045) );
	nand2i_6 U3671 ( .x(n3184), .a(n1657), .b(n3202) );
	nor2i_8 U3672 ( .x(n1174), .a(n634), .b(n1175) );
	inv_16 U3673 ( .x(n3592), .a(n1645) );
	inv_14 U3674 ( .x(n1685), .a(n1624) );
	inv_8 U3675 ( .x(n2070), .a(n1418) );
	inv_16 U3676 ( .x(n1982), .a(n1419) );
	inv_10 U3677 ( .x(n2227), .a(n2128) );
	nand2i_6 U3679 ( .x(n3503), .a(n1577), .b(n927) );
	nand2_2 U368 ( .x(n690), .a(___cell__39620_net147732), .b(___cell__39620_net144201) );
	inv_6 U3680 ( .x(n3517), .a(n3560) );
	nand2i_5 U3683 ( .x(n3567), .a(n1219), .b(n874) );
	nand2i_5 U3685 ( .x(n3361), .a(n1587), .b(n874) );
	nand2i_5 U3686 ( .x(n3297), .a(n1649), .b(n874) );
	nand2i_5 U3687 ( .x(n3363), .a(n1580), .b(n874) );
	nand2i_6 U3689 ( .x(n3372), .a(n1571), .b(n928) );
	oai21_1 U369 ( .x(n3102), .a(n1511), .b(n690), .c(n3103) );
	nand2i_6 U3690 ( .x(n3548), .a(n1572), .b(n927) );
	nand2i_5 U3691 ( .x(n3549), .a(n1646), .b(n874) );
	nand2i_6 U3692 ( .x(n3292), .a(n1529), .b(n928) );
	nand2i_6 U3693 ( .x(n3304), .a(n1570), .b(n928) );
	nand2_8 U3694 ( .x(n3725), .a(___cell__39620_net144328), .b(___cell__39620_net144331) );
	nand2i_6 U3695 ( .x(n3376), .a(n1585), .b(n928) );
	inv_6 U3698 ( .x(n1148), .a(n3394) );
	nand2i_5 U3699 ( .x(n3453), .a(n1579), .b(n874) );
	inv_12 U37 ( .x(n609), .a(n1585) );
	nand2i_0 U370 ( .x(n1388), .a(n1579), .b(n530) );
	nand2_8 U3700 ( .x(n1715), .a(n1691), .b(n1714) );
	nand2i_6 U3701 ( .x(n1713), .a(n1546), .b(n1714) );
	nand2i_6 U3702 ( .x(n3402), .a(n1587), .b(n883) );
	nor2i_5 U3704 ( .x(n1146), .a(n1147), .b(n1148) );
	aoi21_6 U3705 ( .x(n2110), .a(n2066), .b(n686), .c(n2067) );
	inv_10 U3706 ( .x(n2066), .a(n1672) );
	nand2i_6 U3707 ( .x(n1974), .a(n855), .b(n1553) );
	inv_6 U3708 ( .x(n2214), .a(n3340) );
	nand2_8 U3709 ( .x(n1556), .a(n1555), .b(n855) );
	aoi21_1 U371 ( .x(n1387), .a(n1143), .b(n1388), .c(n653) );
	nand2i_6 U3710 ( .x(n3657), .a(n924), .b(n910) );
	nand2i_5 U3711 ( .x(n3574), .a(n924), .b(n901) );
	inv_16 U3712 ( .x(n3575), .a(n4013) );
	nand2i_6 U3713 ( .x(n2115), .a(n1644), .b(n928) );
	nor2_1 U372 ( .x(n1389), .a(n4002), .b(n588) );
	inv_2 U373 ( .x(n1382), .a(N1809) );
	nor2_1 U374 ( .x(n1381), .a(n1077), .b(n1382) );
	inv_12 U375 ( .x(n1579), .a(reg_out_A[12]) );
	ao211_5 U3750 ( .x(n3084), .a(n3110), .b(n1267), .c(n4119), .d(n4118) );
	inv_0 U3751 ( .x(n4118), .a(n3089) );
	inv_2 U3752 ( .x(n4119), .a(n3088) );
	nand2i_1 U3753 ( .x(n3088), .a(n4022), .b(n3057) );
	ao211_5 U3754 ( .x(n2806), .a(n3464), .b(n4122), .c(n4121), .d(n4120) );
	inv_2 U3755 ( .x(n4120), .a(n2216) );
	inv_4 U3756 ( .x(n4121), .a(n3331) );
	inv_0 U3757 ( .x(n4122), .a(___cell__39620_net144317) );
	nand2i_5 U3758 ( .x(n2216), .a(n1649), .b(n4130) );
	nand2_1 U3759 ( .x(n3331), .a(n1686), .b(n749) );
	nor2i_1 U376 ( .x(n1376), .a(n1377), .b(___cell__39620_net143658) );
	ao21_6 U3760 ( .x(n2603), .a(n4124), .b(n3388), .c(n4123) );
	inv_2 U3761 ( .x(n4123), .a(n3461) );
	inv_3 U3762 ( .x(n4124), .a(n4125) );
	inv_14 U3763 ( .x(n4125), .a(___cell__39620_net144317) );
	inv_4 U3764 ( .x(n1152), .a(n3388) );
	nand2i_6 U3765 ( .x(n3388), .a(n3389), .b(n3390) );
	nand3_2 U3766 ( .x(n2868), .a(n730), .b(n2873), .c(n2871) );
	inv_3 U3767 ( .x(___cell__39620_net144317), .a(Imm[3]) );
	inv_12 U3768 ( .x(net149167), .a(n799) );
	nand2i_2 U3769 ( .x(n2897), .a(n1626), .b(n3873) );
	nor2i_1 U377 ( .x(n1378), .a(N1710), .b(___cell__39620_net143660) );
	nand2i_1 U3770 ( .x(n2866), .a(n1641), .b(n3873) );
	oai211_3 U3771 ( .x(n3873), .a(n3529), .b(___cell__39620_net144345), .c(n3871),
		.d(n3872) );
	inv_5 U3772 ( .x(n3130), .a(n2050) );
	aoi21_1 U3773 ( .x(n2049), .a(n1221), .b(n2050), .c(n2046) );
	nand2i_0 U3774 ( .x(n2015), .a(n1588), .b(n2050) );
	oai221_4 U3775 ( .x(n2050), .a(n3439), .b(n1559), .c(n747), .d(n1562),
		.e(n1975) );
	ao222_4 U3776 ( .x(n2908), .a(n2874), .b(n755), .c(n2875), .d(n756), .e(ALU_result[18]),
		.f(n3057) );
	aoi211_2 U3777 ( .x(n730), .a(n2798), .b(n1085), .c(n732), .d(n731) );
	inv_6 U3778 ( .x(n731), .a(n2876) );
	aoi211_1 U3779 ( .x(n998), .a(n977), .b(N348), .c(n2051), .d(n2055) );
	inv_5 U378 ( .x(n3546), .a(n3545) );
	nand2i_3 U3780 ( .x(n3300), .a(n1656), .b(n874) );
	oai21_2 U3781 ( .x(n2898), .a(n1566), .b(n4126), .c(n3890) );
	inv_5 U3782 ( .x(n4126), .a(n2899) );
	nand4i_4 U3783 ( .x(n2899), .a(n1299), .b(n3881), .c(n3880), .d(n3879) );
	inv_16 U3784 ( .x(n649), .a(n1566) );
	nand2i_0 U3785 ( .x(n3890), .a(n1500), .b(n2139) );
	nand2i_5 U3786 ( .x(n1566), .a(___cell__39620_net144175), .b(n1567) );
	nand2_3 U3787 ( .x(n695), .a(n713), .b(n4130) );
	nand2i_2 U3788 ( .x(n2163), .a(n1656), .b(n4130) );
	nand2i_2 U3789 ( .x(n3568), .a(n862), .b(n4130) );
	nor2i_3 U379 ( .x(n1106), .a(___cell__39620_net143722), .b(n746) );
	nand2i_2 U3790 ( .x(n3562), .a(n1648), .b(n4130) );
	nand2i_2 U3791 ( .x(n3364), .a(n748), .b(n4130) );
	nand2i_2 U3792 ( .x(n3686), .a(n1655), .b(n4130) );
	nand2i_2 U3793 ( .x(n3295), .a(n1586), .b(n4130) );
	nand2i_1 U3794 ( .x(n3393), .a(n1587), .b(n4130) );
	oai22_2 U3795 ( .x(n2189), .a(n895), .b(n4001), .c(n3525), .d(n784) );
	aoi211_2 U3796 ( .x(n2879), .a(N1650), .b(n809), .c(n1303), .d(n2878) );
	nor2i_5 U3797 ( .x(n1303), .a(N1716), .b(___cell__39620_net143660) );
	aoi22_2 U3798 ( .x(n2712), .a(n2713), .b(___cell__39620_net143722), .c(___cell__39620_net143864),
		.d(n2714) );
	inv_3 U3799 ( .x(n1205), .a(n2457) );
	nand4_1 U38 ( .x(n3221), .a(n1506), .b(n1504), .c(n1509), .d(n1507) );
	aoi21_1 U380 ( .x(n2084), .a(n1249), .b(n2000), .c(n2082) );
	nand2_1 U3800 ( .x(n4128), .a(n3502), .b(n3503) );
	nand2_2 U3801 ( .x(n4127), .a(n3502), .b(n3503) );
	nand2i_3 U3802 ( .x(n3502), .a(n1578), .b(n874) );
	nand2_1 U3803 ( .x(n3097), .a(n3502), .b(n3503) );
	oai221_1 U3804 ( .x(n4129), .a(n3553), .b(___cell__39620_net144374), .c(n3299),
		.d(n1623), .e(n2853) );
	aoi22_2 U3805 ( .x(n2853), .a(n1066), .b(n2854), .c(n1683), .d(n2563) );
	buf_14 U3806 ( .x(n4130), .a(n531) );
	buf_8 U3807 ( .x(n927), .a(n531) );
	buf_14 U3808 ( .x(n928), .a(n531) );
	nand2_5 U3809 ( .x(n3034), .a(n3359), .b(n3360) );
	nand2_1 U381 ( .x(n3685), .a(n1256), .b(n2187) );
	nand2i_4 U3810 ( .x(n3360), .a(n1569), .b(n928) );
	nand2i_4 U3811 ( .x(n3359), .a(n1573), .b(n874) );
	oai31_2 U3812 ( .x(n1010), .a(n2425), .b(n2413), .c(n2418), .d(___cell__39620_net143326) );
	ao21_6 U3813 ( .x(n3765), .a(n4131), .b(n3723), .c(n4132) );
	inv_0 U3814 ( .x(n4131), .a(net149122) );
	ao22_3 U3815 ( .x(n4132), .a(___cell__39620_net144517), .b(n2279), .c(n1391),
		.d(n2375) );
	buf_16 U3816 ( .x(net149122), .a(net149107) );
	oai211_3 U3817 ( .x(n2302), .a(n550), .b(___cell__39620_net144317), .c(n3392),
		.d(n3393) );
	inv_4 U3818 ( .x(n550), .a(n3496) );
	oai221_2 U3819 ( .x(n3116), .a(n511), .b(n1635), .c(n3335), .d(n4009),
		.e(n3098) );
	aoi21_1 U382 ( .x(n2081), .a(n1714), .b(n1999), .c(n1092) );
	oa22_5 U3820 ( .x(n511), .a(n1570), .b(n1629), .c(n512), .d(n536) );
	inv_7 U3821 ( .x(n912), .a(n911) );
	oai22_1 U3822 ( .x(n4133), .a(n1572), .b(n836), .c(n3397), .d(n4125) );
	oai22_1 U3823 ( .x(n4134), .a(n1572), .b(n836), .c(n3397), .d(n4125) );
	oai22_1 U3824 ( .x(n2563), .a(n1572), .b(n836), .c(n3397), .d(n4125) );
	inv_10 U3825 ( .x(n3397), .a(n3541) );
	nand4_2 U3826 ( .x(n4078), .a(n993), .b(n992), .c(n991), .d(n990) );
	nand4_1 U3827 ( .x(n4077), .a(n1010), .b(n1008), .c(n1009), .d(n1007) );
	aoi22_1 U3828 ( .x(n2739), .a(n1683), .b(n2649), .c(___cell__39620_net144517),
		.d(n4134) );
	nand2i_1 U3829 ( .x(n3829), .a(n1625), .b(n4133) );
	nand2i_2 U383 ( .x(n3679), .a(n1623), .b(n3457) );
	inv_6 U3830 ( .x(n933), .a(n932) );
	inv_10 U3831 ( .x(n934), .a(n932) );
	inv_7 U3832 ( .x(n932), .a(reg_out_A[14]) );
	nand4_2 U3833 ( .x(n2055), .a(n2058), .b(n2057), .c(n579), .d(n2053) );
	nand4_2 U3834 ( .x(n2425), .a(n2422), .b(n2426), .c(n2427), .d(n2424) );
	nand4_3 U3835 ( .x(_ALU_result_reg_31_net106451), .a(___cell__39620_net143598),
		.b(___cell__39620_net143595), .c(___cell__39620_net143597), .d(___cell__39620_net143596) );
	and4i_5 U3836 ( .x(___cell__39620_net143598), .a(n2295), .b(n2299), .c(n2298),
		.d(n2297) );
	nand2i_4 U3837 ( .x(n2426), .a(n1759), .b(n1987) );
	inv_3 U3838 ( .x(n1751), .a(N1859) );
	and4i_3 U3839 ( .x(n990), .a(n2392), .b(n2389), .c(n2404), .d(n2401) );
	nand4_1 U384 ( .x(n3681), .a(n3679), .b(n3678), .c(n3680), .d(n2078) );
	oai211_2 U3840 ( .x(n2392), .a(n2393), .b(n4001), .c(n2394), .d(n2395) );
	aoi211_2 U3841 ( .x(n2073), .a(N1705), .b(___cell__39620_net145190), .c(n1097),
		.d(n1096) );
	aoi22_3 U3842 ( .x(n2385), .a(N1826), .b(n1987), .c(n1095), .d(n2386) );
	inv_14 U3843 ( .x(n637), .a(n738) );
	inv_7 U3844 ( .x(n2429), .a(n2270) );
	nand2_5 U3845 ( .x(n2270), .a(n3563), .b(n3564) );
	inv_4 U3846 ( .x(n931), .a(n929) );
	inv_10 U3847 ( .x(n930), .a(n929) );
	inv_6 U3848 ( .x(n929), .a(reg_out_A[13]) );
	nor2i_2 U3849 ( .x(n1240), .a(N1654), .b(___cell__39620_net143872) );
	nor2_1 U385 ( .x(n1105), .a(___cell__39620_net143693), .b(___cell__39620_net143720) );
	aoai211_4 U3850 ( .x(n4049), .a(___cell__39620_net143287), .b(n1455), .c(n1439),
		.d(n1456) );
	nand2_4 U3851 ( .x(n613), .a(n615), .b(n614) );
	nand2i_2 U3852 ( .x(n3712), .a(n727), .b(n2809) );
	oai211_3 U3853 ( .x(n2809), .a(n3334), .b(n1546), .c(n3339), .d(n3340) );
	nor2_2 U3854 ( .x(n1953), .a(reg_out_B[8]), .b(reg_out_B[9]) );
	nand2i_4 U3855 ( .x(n736), .a(reg_out_B[29]), .b(n1731) );
	inv_0 U3856 ( .x(n4135), .a(net149617) );
	inv_2 U3857 ( .x(n4136), .a(n4135) );
	inv_6 U3858 ( .x(net149617), .a(net149616) );
	nand3_4 U3859 ( .x(n679), .a(n678), .b(n1663), .c(n701) );
	nand2i_2 U386 ( .x(n2087), .a(n1461), .b(n2139) );
	inv_6 U3860 ( .x(n701), .a(___cell__39620_net144175) );
	buf_2 U3861 ( .x(n4015), .a(reg_out_A[1]) );
	and2_1 U3862 ( .x(n4137), .a(n4138), .b(IR_opcode_field[4]) );
	inv_2 U3863 ( .x(n1609), .a(n4137) );
	inv_0 U3864 ( .x(n4138), .a(IR_opcode_field[5]) );
	buf_8 U3865 ( .x(net149107), .a(Imm[1]) );
	inv_10 U3866 ( .x(n896), .a(n1554) );
	nand2i_8 U3867 ( .x(n1554), .a(reg_out_B[5]), .b(n1552) );
	and2_5 U3868 ( .x(n1241), .a(N1720), .b(___cell__39620_net145190) );
	nand2i_4 U3869 ( .x(___cell__39620_net143660), .a(IR_opcode_field[2]),
		.b(___cell__39620_net144309) );
	inv_2 U387 ( .x(n3688), .a(n1462) );
	inv_16 U3870 ( .x(___cell__39620_net145190), .a(___cell__39620_net143660) );
	nand2i_2 U3871 ( .x(n2152), .a(n1641), .b(n3689) );
	nand2i_2 U3872 ( .x(n2257), .a(n1641), .b(n3711) );
	nand2i_4 U3873 ( .x(n2895), .a(n1641), .b(n3887) );
	nand2i_2 U3874 ( .x(n2407), .a(n1641), .b(n2455) );
	nand2i_2 U3875 ( .x(n2976), .a(n1641), .b(n3009) );
	nand2i_1 U3876 ( .x(n2029), .a(n1641), .b(n3583) );
	nand2i_2 U3877 ( .x(n2102), .a(n1641), .b(n3681) );
	oai22_2 U3878 ( .x(n2489), .a(n621), .b(n1122), .c(n1641), .d(n1120) );
	nand2i_2 U3879 ( .x(n3143), .a(n1641), .b(n3168) );
	nand2_2 U388 ( .x(n2086), .a(n2193), .b(n3688) );
	inv_3 U3880 ( .x(n905), .a(Imm[13]) );
	inv_2 U3881 ( .x(n555), .a(Imm[13]) );
	aoi22_3 U3882 ( .x(n2312), .a(N1827), .b(n1987), .c(N1860), .d(n4000) );
	nand2_2 U3883 ( .x(n1632), .a(n816), .b(reg_out_B[2]) );
	or2_6 U3884 ( .x(n1565), .a(reg_out_B[2]), .b(reg_out_B[3]) );
	nand2_1 U3885 ( .x(n1634), .a(n879), .b(reg_out_B[2]) );
	inv_7 U3886 ( .x(n828), .a(reg_out_B[2]) );
	buf_10 U3887 ( .x(n608), .a(reg_out_A[15]) );
	buf_4 U3888 ( .x(n4139), .a(reg_out_B[21]) );
	buf_8 U3889 ( .x(n918), .a(n931) );
	oai211_1 U389 ( .x(n2085), .a(n1104), .b(n1671), .c(n2086), .d(n2087) );
	buf_6 U3890 ( .x(n4014), .a(reg_out_A[15]) );
	buf_5 U3891 ( .x(n4016), .a(reg_out_A[15]) );
	buf_4 U3892 ( .x(n602), .a(reg_out_A[15]) );
	nand2_8 U3893 ( .x(n4140), .a(___cell__39620_net144330), .b(reg_out_A[31]) );
	inv_10 U3894 ( .x(n817), .a(Imm[10]) );
	or3i_5 U3895 ( .x(n1957), .a(n605), .b(reg_out_B[20]), .c(reg_out_B[18]) );
	nand4i_1 U3896 ( .x(n4141), .a(n1360), .b(n3968), .c(n3967), .d(n3966) );
	oai211_2 U3897 ( .x(n4069), .a(n1020), .b(___cell__39620_net143287), .c(n1021),
		.d(n1022) );
	ao21_4 U3898 ( .x(n4142), .a(net150830), .b(n2080), .c(n837) );
	inv_5 U3899 ( .x(n837), .a(n3456) );
	exnor2_1 U39 ( .x(n3231), .a(net152465), .b(n942) );
	nor2_1 U390 ( .x(n1107), .a(n1087), .b(n4043) );
	ao211_2 U3900 ( .x(n4067), .a(___cell__39620_net143326), .b(n974), .c(n975),
		.d(n976) );
	nand4i_2 U3901 ( .x(n974), .a(n1309), .b(n2882), .c(n2881), .d(n2883) );
	inv_16 U3902 ( .x(N69), .a(reg_out_A[31]) );
	nand2_8 U3903 ( .x(n1159), .a(n896), .b(reg_out_A[31]) );
	inv_0 U3904 ( .x(n4143), .a(reg_out_B[31]) );
	inv_2 U3905 ( .x(n4144), .a(n4143) );
	nor2_2 U3906 ( .x(n1955), .a(reg_out_B[13]), .b(reg_out_B[14]) );
	inv_6 U3907 ( .x(n4145), .a(reg_out_B[7]) );
	inv_10 U3908 ( .x(n4146), .a(n4145) );
	inv_5 U3909 ( .x(n759), .a(reg_out_B[5]) );
	oai22_2 U391 ( .x(n2135), .a(n890), .b(n1656), .c(n1651), .d(n1657) );
	buf_1 U3910 ( .x(n4147), .a(reg_out_B[9]) );
	buf_16 U3911 ( .x(mem_to_reg_EX), .a(n4224) );
	nor2_1 U3912 ( .x(n1952), .a(reg_out_B[6]), .b(n4146) );
	nor2_2 U3913 ( .x(n1958), .a(reg_out_B[23]), .b(reg_out_B[24]) );
	nor2_3 U3914 ( .x(n1959), .a(reg_out_B[25]), .b(reg_out_B[26]) );
	nor2_1 U3915 ( .x(n1954), .a(reg_out_B[10]), .b(reg_out_B[11]) );
	nor2i_0 U3916 ( .x(n4156), .a(reg_out_B[24]), .b(n4116) );
	and2_1 U3917 ( .x(n4158), .a(reg_out_B[15]), .b(n4117) );
	nor2i_0 U3918 ( .x(n4160), .a(n816), .b(___cell__6067_net21981) );
	nor2i_0 U3919 ( .x(n4162), .a(n566), .b(n4116) );
	inv_5 U392 ( .x(n852), .a(n851) );
	nor2i_0 U3920 ( .x(n4164), .a(reg_out_B[30]), .b(n4116) );
	nor2i_0 U3921 ( .x(n4166), .a(reg_out_B[28]), .b(n4116) );
	nor2i_0 U3922 ( .x(n4168), .a(reg_out_B[27]), .b(n4116) );
	nor2i_0 U3923 ( .x(n4170), .a(reg_out_B[25]), .b(n4116) );
	nor2i_0 U3924 ( .x(n4172), .a(reg_out_B[23]), .b(n4116) );
	nor2i_0 U3925 ( .x(n4174), .a(reg_out_B[19]), .b(n4116) );
	nor2i_0 U3926 ( .x(n4176), .a(reg_out_B[16]), .b(n4116) );
	and2_1 U3927 ( .x(n4178), .a(reg_out_B[14]), .b(n4117) );
	and2_1 U3928 ( .x(n4180), .a(reg_out_B[12]), .b(n4117) );
	and2_1 U3929 ( .x(n4182), .a(reg_out_B[10]), .b(n4117) );
	inv_2 U393 ( .x(n3793), .a(n1479) );
	and2_1 U3930 ( .x(n4184), .a(reg_out_B[8]), .b(n4117) );
	nor2i_0 U3931 ( .x(n4186), .a(n4146), .b(___cell__6067_net21981) );
	nor2i_0 U3932 ( .x(n4188), .a(reg_out_B[6]), .b(___cell__6067_net21981) );
	nor2i_0 U3933 ( .x(n4190), .a(reg_out_B[5]), .b(___cell__6067_net21981) );
	nor2i_0 U3934 ( .x(n4192), .a(reg_out_B[4]), .b(___cell__6067_net21981) );
	nor2i_0 U3935 ( .x(n4194), .a(n536), .b(___cell__6067_net21981) );
	nor2i_0 U3936 ( .x(n4196), .a(n815), .b(___cell__6067_net21981) );
	and2_1 U3937 ( .x(n4198), .a(reg_write), .b(N3304) );
	and2_1 U3938 ( .x(n4200), .a(mem_to_reg), .b(N3304) );
	and2_1 U3939 ( .x(n4202), .a(mem_read), .b(N3304) );
	nand2_2 U394 ( .x(n2483), .a(n2193), .b(n3793) );
	and2_1 U3940 ( .x(n4203), .a(mem_write), .b(N3304) );
	nor2i_0 U3941 ( .x(n4204), .a(reg_out_B[22]), .b(n4116) );
	nor2i_0 U3942 ( .x(n4206), .a(reg_out_B[26]), .b(n4116) );
	and2_1 U3943 ( .x(n4208), .a(n4147), .b(n4117) );
	nor2i_0 U3944 ( .x(n4210), .a(reg_out_B[18]), .b(n4116) );
	nor2i_0 U3945 ( .x(n4212), .a(reg_out_B[0]), .b(___cell__6067_net21981) );
	and2_1 U3946 ( .x(n4214), .a(reg_out_B[11]), .b(n4117) );
	and2_1 U3947 ( .x(n4216), .a(reg_out_B[13]), .b(n4117) );
	nor2i_0 U3948 ( .x(n4218), .a(reg_out_B[20]), .b(n4116) );
	nor2i_0 U3949 ( .x(n4220), .a(reg_out_B[29]), .b(n4116) );
	nand2i_2 U395 ( .x(n2482), .a(n1480), .b(n2139) );
	nor2i_0 U3950 ( .x(n4222), .a(reg_out_B[17]), .b(n4116) );
	oa22_2 U396 ( .x(n505), .a(n1637), .b(n1093), .c(n1626), .d(n1089) );
	oai211_1 U397 ( .x(n2481), .a(n505), .b(n1580), .c(n2482), .d(n2483) );
	nand2i_3 U398 ( .x(n2487), .a(n2459), .b(n866) );
	inv_2 U399 ( .x(n3792), .a(n3791) );
	nand4_1 U40 ( .x(n3230), .a(n3231), .b(n1458), .c(n1462), .d(n1460) );
	nand2i_2 U400 ( .x(n2461), .a(n816), .b(n502) );
	nand2i_2 U401 ( .x(n2485), .a(n2461), .b(n3778) );
	nand2_2 U402 ( .x(n3743), .a(n3477), .b(___cell__39620_net144331) );
	inv_2 U403 ( .x(n1766), .a(N1758) );
	nand2i_2 U404 ( .x(n2468), .a(n1766), .b(___cell__39620_net145150) );
	nand2i_0 U405 ( .x(n2467), .a(___cell__39620_net144655), .b(n663) );
	nand2_2 U406 ( .x(n2462), .a(n681), .b(n537) );
	nand2i_2 U407 ( .x(n2464), .a(n2462), .b(___cell__39620_net145285) );
	inv_2 U408 ( .x(n1933), .a(N1797) );
	inv_2 U409 ( .x(n1936), .a(N1830) );
	inv_2 U41 ( .x(n2194), .a(n1465) );
	oai22_1 U410 ( .x(n3252), .a(n946), .b(n1936), .c(n1077), .d(n1933) );
	inv_2 U411 ( .x(n1930), .a(N1731) );
	inv_2 U412 ( .x(n1929), .a(N1698) );
	oai221_1 U413 ( .x(n3249), .a(___cell__39620_net143660), .b(n1929), .c(___cell__39620_net143710),
		.d(n1930), .e(n3250) );
	ao211_3 U414 ( .x(n3251), .a(n1318), .b(n1423), .c(n3249), .d(n3252) );
	nand2i_2 U415 ( .x(n3255), .a(n1934), .b(n3624) );
	inv_2 U416 ( .x(n1934), .a(N1996) );
	inv_2 U417 ( .x(n1932), .a(N1930) );
	nand2i_2 U418 ( .x(n3254), .a(n1932), .b(n3662) );
	nand2i_2 U419 ( .x(n3253), .a(n1935), .b(___cell__39620_net145508) );
	inv_5 U42 ( .x(net152465), .a(n783) );
	inv_2 U420 ( .x(n1935), .a(N1963) );
	nor2i_1 U421 ( .x(n1438), .a(N1632), .b(___cell__39620_net143872) );
	nor2i_3 U422 ( .x(n1435), .a(n1436), .b(n1437) );
	aoi21_1 U423 ( .x(n3240), .a(net152465), .b(n3241), .c(n701) );
	aoai211_1 U424 ( .x(n3243), .a(n891), .b(n3539), .c(n3236), .d(n1095) );
	oai211_2 U425 ( .x(n3242), .a(n1430), .b(n1639), .c(n3243), .d(n3240) );
	oai21_1 U426 ( .x(n3237), .a(n1427), .b(n1089), .c(n1618) );
	inv_1 U427 ( .x(n545), .a(n889) );
	exnor2_1 U428 ( .x(n1945), .a(n3990), .b(___cell__39620_net144166) );
	ao222_2 U429 ( .x(n742), .a(n1256), .b(n2809), .c(n2273), .d(n893), .e(n1150),
		.f(n3279) );
	nand2i_0 U43 ( .x(n1527), .a(n1524), .b(n1528) );
	inv_5 U430 ( .x(n3860), .a(n1836) );
	inv_2 U431 ( .x(n1567), .a(n1544) );
	aoai211_1 U432 ( .x(n3286), .a(n3591), .b(n1567), .c(n3280), .d(n942) );
	nand2i_2 U433 ( .x(n1544), .a(n816), .b(n1545) );
	nand2i_2 U434 ( .x(n3285), .a(n1560), .b(n3715) );
	aoi21_1 U435 ( .x(n3277), .a(n1177), .b(n3278), .c(n3276) );
	aoai211_1 U436 ( .x(n3284), .a(n3277), .b(n3285), .c(n1544), .d(n3286) );
	exnor2_1 U437 ( .x(n1949), .a(n1950), .b(n1530) );
	mux2i_2 U438 ( .x(n3994), .d0(n1947), .sl(IR_function_field[0]), .d1(N1402) );
	oaoi211_1 U439 ( .x(n1445), .a(n942), .b(n1446), .c(n1447), .d(n1448) );
	nand4_1 U44 ( .x(n3259), .a(n1505), .b(n1503), .c(n1510), .d(n1508) );
	nand2i_2 U440 ( .x(n1447), .a(n1531), .b(n1528) );
	inv_1 U441 ( .x(n1448), .a(reg_out_B[0]) );
	inv_2 U442 ( .x(n1537), .a(n1446) );
	nor2i_1 U443 ( .x(n1453), .a(N307), .b(n1454) );
	inv_2 U444 ( .x(n1593), .a(n1454) );
	nand2i_2 U445 ( .x(n3128), .a(n1513), .b(n2139) );
	exnor2_1 U446 ( .x(n1514), .a(n753), .b(n901) );
	inv_2 U447 ( .x(n3982), .a(n1514) );
	nand2_2 U448 ( .x(n3127), .a(n2193), .b(n3982) );
	aoi21_1 U449 ( .x(n1403), .a(n901), .b(n530), .c(n1064) );
	inv_0 U45 ( .x(n1916), .a(reg_out_B[10]) );
	inv_4 U450 ( .x(n1300), .a(n3022) );
	inv_3 U451 ( .x(n3417), .a(n3415) );
	nor2_0 U452 ( .x(n1404), .a(n1087), .b(n4021) );
	ao22_2 U453 ( .x(n716), .a(n1391), .b(n3034), .c(n1066), .d(n3097) );
	ao221_4 U454 ( .x(n3113), .a(n3451), .b(n715), .c(n714), .d(n713), .e(n716) );
	nor2i_1 U455 ( .x(n1398), .a(N1841), .b(n946) );
	nor2i_0 U456 ( .x(n1394), .a(n753), .b(n1586) );
	nor2i_0 U457 ( .x(n1393), .a(n1394), .b(___cell__39620_net143658) );
	nor2i_3 U458 ( .x(n1395), .a(N1709), .b(___cell__39620_net143660) );
	inv_2 U459 ( .x(n1912), .a(N1874) );
	nand3_1 U46 ( .x(n3258), .a(n1513), .b(n1512), .c(n1515) );
	inv_5 U460 ( .x(n3459), .a(n2262) );
	nor2_1 U461 ( .x(n1269), .a(n679), .b(n4027) );
	exnor2_1 U462 ( .x(n1494), .a(n749), .b(n551) );
	inv_2 U463 ( .x(n2787), .a(n1494) );
	inv_2 U464 ( .x(n2786), .a(n1493) );
	aoi22_1 U465 ( .x(n2785), .a(n2139), .b(n2786), .c(n2193), .d(n2787) );
	inv_2 U466 ( .x(n1259), .a(n3020) );
	ao22_2 U467 ( .x(n2772), .a(n661), .b(n662), .c(net151904), .d(n663) );
	inv_2 U468 ( .x(n1826), .a(N1652) );
	nand2i_2 U469 ( .x(n2771), .a(n1826), .b(n809) );
	inv_0 U47 ( .x(n1771), .a(reg_out_B[26]) );
	nand2_2 U470 ( .x(n2764), .a(n551), .b(n749) );
	nand2i_2 U471 ( .x(n2770), .a(n2764), .b(___cell__39620_net147791) );
	inv_5 U472 ( .x(n3656), .a(n3655) );
	nand2i_2 U473 ( .x(n3043), .a(n1508), .b(n2139) );
	oai21_1 U474 ( .x(n3042), .a(n1507), .b(n690), .c(n3043) );
	nand2i_2 U475 ( .x(n1357), .a(n1571), .b(n530) );
	aoi21_1 U476 ( .x(n1356), .a(n1143), .b(n1357), .c(n1358) );
	nor2_1 U477 ( .x(n1359), .a(n4002), .b(___cell__39620_net143997) );
	nand2i_2 U478 ( .x(n3964), .a(n703), .b(n3013) );
	nor2_1 U48 ( .x(n3268), .a(n3269), .b(n3270) );
	inv_2 U480 ( .x(n1887), .a(N1877) );
	nand2i_2 U481 ( .x(n3027), .a(n1887), .b(n944) );
	nand2i_2 U482 ( .x(n3026), .a(n3023), .b(___cell__39620_net147791) );
	nand2i_2 U483 ( .x(n3025), .a(n1886), .b(n809) );
	inv_2 U484 ( .x(n1886), .a(N1646) );
	nor2i_1 U485 ( .x(n1350), .a(N1712), .b(___cell__39620_net143660) );
	nand2i_2 U486 ( .x(n3937), .a(n1043), .b(n3538) );
	nor2i_3 U487 ( .x(n1323), .a(n1147), .b(n1324) );
	nand2i_2 U488 ( .x(n3973), .a(n1510), .b(n2139) );
	inv_2 U489 ( .x(n1373), .a(n1509) );
	nor2_1 U49 ( .x(n3265), .a(n3266), .b(n3267) );
	nor2i_1 U490 ( .x(n1372), .a(n1373), .b(n690) );
	nand2i_2 U491 ( .x(n3970), .a(n727), .b(n2852) );
	nand2_2 U493 ( .x(n702), .a(n701), .b(n1661) );
	nand2i_2 U494 ( .x(n1370), .a(n1563), .b(n530) );
	aoi21_1 U495 ( .x(n1369), .a(n1143), .b(n1370), .c(n1371) );
	oa22_2 U499 ( .x(n849), .a(n3345), .b(n536), .c(n1561), .d(n1629) );
	inv_2 U50 ( .x(n2195), .a(n1466) );
	nand2i_2 U500 ( .x(n3965), .a(___cell__39620_net144062), .b(n3457) );
	aoi21_4 U501 ( .x(n630), .a(net150830), .b(n2080), .c(n837) );
	nand2i_0 U502 ( .x(n3089), .a(n1563), .b(n1700) );
	nor2_1 U504 ( .x(n1374), .a(___cell__39620_net143693), .b(n1375) );
	aoi22_1 U505 ( .x(n3032), .a(n1391), .b(n3033), .c(n1066), .d(n3034) );
	nand2i_2 U506 ( .x(n3957), .a(___cell__39620_net144374), .b(n4128) );
	inv_0 U507 ( .x(n1371), .a(reg_out_B[13]) );
	nor2i_1 U508 ( .x(n1364), .a(N1843), .b(n946) );
	inv_2 U509 ( .x(n1895), .a(N1876) );
	inv_8 U51 ( .x(n682), .a(___cell__39620_net144029) );
	nand2i_2 U510 ( .x(n3063), .a(n1895), .b(n3998) );
	nor2i_1 U511 ( .x(n1362), .a(N1711), .b(___cell__39620_net143660) );
	inv_14 U512 ( .x(n708), .a(___cell__39620_net144170) );
	inv_2 U513 ( .x(___cell__39620_net145285), .a(___cell__39620_net143658) );
	aoi21_1 U515 ( .x(n3061), .a(n3060), .b(___cell__39620_net145285), .c(n1362) );
	inv_2 U516 ( .x(n3157), .a(n1516) );
	exnor2_1 U517 ( .x(n1515), .a(n908), .b(reg_out_B[10]) );
	inv_2 U518 ( .x(n3156), .a(n1515) );
	aoi22_1 U519 ( .x(n3155), .a(n2139), .b(n3156), .c(n2193), .d(n3157) );
	nand2i_2 U520 ( .x(n3159), .a(n1916), .b(n530) );
	inv_5 U521 ( .x(n1313), .a(n3059) );
	inv_8 U522 ( .x(n3358), .a(n3356) );
	oai22_3 U523 ( .x(n3516), .a(n1649), .b(n1651), .c(n3517), .d(n891) );
	inv_2 U524 ( .x(n3513), .a(n3863) );
	nand2i_2 U525 ( .x(n3512), .a(n3513), .b(n3514) );
	inv_5 U526 ( .x(n3413), .a(n3410) );
	oai22_1 U527 ( .x(n850), .a(n915), .b(n1649), .c(n508), .d(n815) );
	inv_5 U528 ( .x(n3411), .a(n3544) );
	nor2_1 U529 ( .x(n1415), .a(n1087), .b(n4020) );
	nor2_5 U53 ( .x(n775), .a(Imm[18]), .b(Imm[21]) );
	nor2i_2 U530 ( .x(n1414), .a(n502), .b(n720) );
	nand2i_2 U531 ( .x(n3975), .a(n719), .b(n3457) );
	inv_2 U532 ( .x(n1392), .a(n2991) );
	nand4_1 U533 ( .x(n3981), .a(n3980), .b(n3979), .c(n3978), .d(n3977) );
	nand2i_2 U534 ( .x(n3978), .a(n1634), .b(n521) );
	inv_2 U535 ( .x(n3140), .a(n3981) );
	nor2i_1 U536 ( .x(n1409), .a(N1840), .b(n946) );
	nand2i_2 U537 ( .x(n3968), .a(n1608), .b(n3638) );
	nand4i_1 U538 ( .x(n1397), .a(n1360), .b(n3968), .c(n3967), .d(n3966) );
	nor2i_1 U539 ( .x(n1408), .a(N1741), .b(___cell__39620_net143710) );
	inv_3 U54 ( .x(n780), .a(Imm[6]) );
	nor2i_1 U540 ( .x(n1405), .a(n1406), .b(___cell__39620_net143658) );
	nor2i_1 U541 ( .x(n1407), .a(N1708), .b(___cell__39620_net143660) );
	inv_2 U542 ( .x(n3848), .a(n3847) );
	nand2i_2 U543 ( .x(n3847), .a(n601), .b(n530) );
	exnor2_1 U544 ( .x(n1490), .a(n583), .b(n745) );
	inv_2 U545 ( .x(n2694), .a(n1490) );
	exnor2_1 U546 ( .x(n1489), .a(n583), .b(reg_out_B[22]) );
	inv_2 U547 ( .x(n2693), .a(n1489) );
	aoi22_1 U548 ( .x(n2692), .a(n2139), .b(n2693), .c(n2193), .d(n2694) );
	nand2i_2 U549 ( .x(n3849), .a(n601), .b(n1064) );
	nor2_1 U55 ( .x(___cell__39620_net145078), .a(Imm[9]), .b(Imm[15]) );
	nand2i_2 U550 ( .x(n2681), .a(___cell__39620_net143735), .b(n663) );
	inv_2 U551 ( .x(n663), .a(n734) );
	inv_2 U552 ( .x(n1811), .a(N1753) );
	nand2i_2 U553 ( .x(n2680), .a(n1811), .b(___cell__39620_net145150) );
	inv_5 U554 ( .x(n3421), .a(n3774) );
	inv_5 U555 ( .x(n1324), .a(n2766) );
	nand2i_2 U556 ( .x(n2679), .a(n1055), .b(n2600) );
	nor2i_0 U558 ( .x(n2674), .a(n745), .b(n1570) );
	nand2_2 U559 ( .x(n3818), .a(n3480), .b(___cell__39620_net144331) );
	nor2_0 U56 ( .x(n1979), .a(Imm[22]), .b(Imm[23]) );
	aoi21_1 U560 ( .x(n1130), .a(n1131), .b(n1132), .c(n816) );
	nand2i_2 U561 ( .x(n1131), .a(n702), .b(n2136) );
	nand2i_2 U562 ( .x(n1132), .a(___cell__39620_net144406), .b(n750) );
	nand2i_2 U563 ( .x(n3708), .a(n759), .b(n530) );
	inv_2 U564 ( .x(n3709), .a(n3708) );
	exnor2_1 U565 ( .x(n1466), .a(n912), .b(reg_out_B[5]) );
	nand2i_2 U566 ( .x(n2210), .a(n4041), .b(n3057) );
	oai211_2 U567 ( .x(n3689), .a(n3505), .b(n718), .c(n2126), .d(n2127) );
	oai22_1 U568 ( .x(n2205), .a(___cell__39620_net144326), .b(n4002), .c(n2206),
		.d(n1654) );
	inv_2 U569 ( .x(n2366), .a(n2148) );
	nor2_1 U57 ( .x(n1980), .a(Imm[25]), .b(Imm[27]) );
	nand2i_2 U570 ( .x(n2204), .a(n1646), .b(n2148) );
	nand2i_2 U571 ( .x(n2203), .a(n759), .b(n1064) );
	aoi21_1 U572 ( .x(n2132), .a(n1249), .b(n2133), .c(n2131) );
	aoi21_1 U573 ( .x(n2129), .a(n1714), .b(n2130), .c(n1110) );
	nand3_1 U574 ( .x(n3693), .a(n2129), .b(n3692), .c(n2132) );
	inv_5 U575 ( .x(net151578), .a(net151577) );
	inv_2 U576 ( .x(n1125), .a(N1868) );
	nor2_1 U577 ( .x(n1124), .a(n947), .b(n1125) );
	nor2i_3 U578 ( .x(n1297), .a(n650), .b(n1298) );
	inv_2 U579 ( .x(n2630), .a(n3570) );
	inv_2 U58 ( .x(n688), .a(Imm[25]) );
	oai211_1 U580 ( .x(n743), .a(n3600), .b(n1565), .c(n3845), .d(n2672) );
	nand2i_2 U581 ( .x(n3874), .a(n1843), .b(n530) );
	inv_2 U582 ( .x(n3875), .a(n3874) );
	nand2i_2 U583 ( .x(n2870), .a(n1843), .b(n1064) );
	oai21_1 U584 ( .x(n2869), .a(___cell__39620_net143693), .b(n683), .c(n2870) );
	inv_4 U585 ( .x(n1268), .a(n2872) );
	nand2i_2 U586 ( .x(n3519), .a(n3520), .b(n3521) );
	and2_1 U588 ( .x(n732), .a(ALU_result[19]), .b(n3057) );
	inv_2 U589 ( .x(n1292), .a(N1816) );
	nand2i_3 U59 ( .x(n1729), .a(n1043), .b(n1685) );
	nor2_1 U590 ( .x(n1291), .a(n1077), .b(n1292) );
	inv_2 U592 ( .x(n1846), .a(N1717) );
	nand2i_2 U593 ( .x(n2844), .a(n1846), .b(___cell__39620_net145190) );
	nor2i_0 U594 ( .x(n2839), .a(n684), .b(n1583) );
	inv_2 U595 ( .x(n1847), .a(N1750) );
	nand2i_2 U596 ( .x(n3440), .a(n4003), .b(n1977) );
	nand2i_3 U597 ( .x(n3606), .a(n3605), .b(n3598) );
	inv_5 U598 ( .x(n3442), .a(n2236) );
	nand2i_0 U599 ( .x(n1144), .a(n1649), .b(n530) );
	inv_2 U60 ( .x(n3573), .a(n1729) );
	aoi21_1 U600 ( .x(n1142), .a(n1143), .b(n1144), .c(n855) );
	nor2i_1 U601 ( .x(n2212), .a(n1085), .b(n816) );
	nor2i_1 U602 ( .x(n2211), .a(___cell__39620_net144345), .b(n1658) );
	exnor2_1 U603 ( .x(n1468), .a(reg_out_B[4]), .b(n834) );
	exnor2_1 U604 ( .x(n1467), .a(n834), .b(net151904) );
	nor2_1 U605 ( .x(n1145), .a(n679), .b(n4040) );
	nand2i_2 U606 ( .x(n2255), .a(n621), .b(n2371) );
	nand2i_2 U607 ( .x(n2252), .a(n1646), .b(n3705) );
	nand2i_2 U608 ( .x(n2251), .a(n1657), .b(n2148) );
	inv_5 U609 ( .x(___cell__39620_net145617), .a(___cell__39620_net143693) );
	nand2_2 U61 ( .x(n1835), .a(n3573), .b(n910) );
	nand2_0 U610 ( .x(n2249), .a(___cell__39620_net145617), .b(net151904) );
	nand3_2 U611 ( .x(n2247), .a(n2180), .b(n3700), .c(n2178) );
	nand2i_2 U612 ( .x(n3700), .a(___cell__39620_net144062), .b(n2337) );
	nor2i_1 U613 ( .x(n1137), .a(N1702), .b(___cell__39620_net143660) );
	nand2i_2 U614 ( .x(n3507), .a(n4006), .b(n1049) );
	nor2i_0 U615 ( .x(n2215), .a(net151904), .b(n1649) );
	inv_5 U616 ( .x(n1649), .a(n834) );
	inv_2 U617 ( .x(n672), .a(n1047) );
	oai211_2 U618 ( .x(n3687), .a(n1334), .b(___cell__39620_net144317), .c(n2069),
		.d(n3686) );
	inv_5 U619 ( .x(n3510), .a(n3687) );
	nand2_0 U62 ( .x(n3630), .a(___cell__39620_net144330), .b(n541) );
	nor2i_1 U620 ( .x(n1123), .a(n1045), .b(n4006) );
	inv_12 U621 ( .x(n1607), .a(n673) );
	inv_8 U622 ( .x(n885), .a(n1654) );
	inv_12 U623 ( .x(n586), .a(n1417) );
	inv_2 U625 ( .x(n3299), .a(n2927) );
	ao22_1 U626 ( .x(n3552), .a(reg_out_A[8]), .b(n3575), .c(n2277), .d(n799) );
	oai221_2 U627 ( .x(n2875), .a(n3553), .b(___cell__39620_net144374), .c(n3299),
		.d(n1623), .e(n2853) );
	aoi23_1 U628 ( .x(n2850), .a(n1249), .b(n2852), .c(n879), .d(n2851), .e(reg_out_B[2]) );
	inv_5 U629 ( .x(n3522), .a(n3519) );
	nand2i_2 U63 ( .x(n1673), .a(reg_out_B[3]), .b(reg_out_B[4]) );
	nand2i_2 U630 ( .x(n2894), .a(n621), .b(n2930) );
	exnor2_1 U631 ( .x(n1499), .a(n910), .b(n633) );
	inv_2 U632 ( .x(n1311), .a(n1499) );
	nor2i_1 U633 ( .x(n1310), .a(n1311), .b(n690) );
	oai21_1 U636 ( .x(n3374), .a(n815), .b(n528), .c(n3375) );
	and2_1 U637 ( .x(n697), .a(n767), .b(n3381) );
	inv_4 U638 ( .x(n3381), .a(n853) );
	inv_2 U639 ( .x(n3889), .a(n3888) );
	nand2i_1 U64 ( .x(n3449), .a(n1219), .b(n1689) );
	inv_2 U640 ( .x(n1854), .a(N1948) );
	inv_2 U641 ( .x(n1855), .a(N1815) );
	nand2i_2 U642 ( .x(n3859), .a(n1608), .b(n3774) );
	inv_2 U643 ( .x(n2634), .a(n3569) );
	aoi21_2 U644 ( .x(n2765), .a(n2676), .b(n2766), .c(n2634) );
	nand2_2 U645 ( .x(n2877), .a(n633), .b(n910) );
	oai22_1 U646 ( .x(n2878), .a(n1602), .b(n734), .c(___cell__39620_net143658),
		.d(n2877) );
	inv_4 U648 ( .x(n1306), .a(N1881) );
	nand2i_2 U649 ( .x(n3869), .a(n1608), .b(n3790) );
	nand2_0 U65 ( .x(n3635), .a(___cell__39620_net144330), .b(n590) );
	nand2i_4 U650 ( .x(n2310), .a(n1734), .b(___cell__39620_net145508) );
	inv_4 U651 ( .x(n1734), .a(N1993) );
	nand2_2 U652 ( .x(n2307), .a(Imm[30]), .b(n535) );
	nand2i_2 U653 ( .x(n2309), .a(n2307), .b(___cell__39620_net147791) );
	inv_2 U654 ( .x(n1735), .a(N1960) );
	nand2i_2 U655 ( .x(n2311), .a(n1735), .b(n3999) );
	nor2i_1 U656 ( .x(n1161), .a(n1095), .b(n1162) );
	inv_8 U657 ( .x(n3524), .a(n3744) );
	nand2i_2 U658 ( .x(n2316), .a(n1737), .b(n3624) );
	inv_2 U659 ( .x(n1737), .a(N2026) );
	nand2_0 U66 ( .x(n3653), .a(___cell__39620_net144330), .b(n540) );
	nand2i_0 U661 ( .x(n3749), .a(n1731), .b(n1064) );
	inv_10 U662 ( .x(n1731), .a(reg_out_B[30]) );
	ao221_4 U663 ( .x(n1733), .a(n737), .b(n597), .c(n598), .d(n599), .e(n1700) );
	nand2i_0 U664 ( .x(n3747), .a(n1731), .b(n530) );
	nand3i_1 U665 ( .x(n2318), .a(n1732), .b(n3747), .c(n3216) );
	inv_2 U666 ( .x(n3748), .a(n1471) );
	nand2_2 U667 ( .x(n2321), .a(n2193), .b(n3748) );
	oai211_1 U668 ( .x(n2320), .a(n578), .b(n1566), .c(n2321), .d(n2322) );
	nand2i_0 U669 ( .x(n2300), .a(___cell__39620_net144175), .b(n1576) );
	inv_10 U67 ( .x(___cell__39620_net144330), .a(___cell__39620_net144329) );
	inv_5 U670 ( .x(n1576), .a(n1160) );
	inv_2 U671 ( .x(n725), .a(n815) );
	nor2i_1 U672 ( .x(___cell__39620_net145451), .a(n504), .b(n670) );
	inv_12 U673 ( .x(n1587), .a(reg_out_A[27]) );
	exnor2_1 U674 ( .x(n1477), .a(reg_out_A[28]), .b(Imm[28]) );
	exnor2_1 U675 ( .x(n1478), .a(reg_out_A[28]), .b(reg_out_B[28]) );
	inv_2 U676 ( .x(n3267), .a(n1478) );
	nor2i_5 U677 ( .x(n1190), .a(n1191), .b(n578) );
	inv_2 U678 ( .x(n2411), .a(n3775) );
	oai22_1 U679 ( .x(n1732), .a(n621), .b(n1093), .c(n1641), .d(n1089) );
	inv_2 U68 ( .x(n1647), .a(n942) );
	nand2i_2 U680 ( .x(n2448), .a(___cell__39620_net144257), .b(n2489) );
	inv_5 U681 ( .x(n3419), .a(n2719) );
	nand2i_2 U682 ( .x(n2447), .a(n1574), .b(n2399) );
	oai21_3 U683 ( .x(n2492), .a(n3418), .b(n1565), .c(n3571) );
	nor2_1 U684 ( .x(n1192), .a(n679), .b(n4035) );
	nand4_1 U685 ( .x(n2457), .a(n2437), .b(n3771), .c(n2434), .d(n3770) );
	nand2i_2 U686 ( .x(n3771), .a(___cell__39620_net144062), .b(n2302) );
	aoi22_1 U687 ( .x(n2434), .a(n2435), .b(n2262), .c(n2436), .d(n904) );
	aoi21_1 U688 ( .x(n2430), .a(n1256), .b(n2306), .c(n2428) );
	nand2i_2 U689 ( .x(n3769), .a(n1636), .b(n2305) );
	nand2i_2 U69 ( .x(n3561), .a(n1647), .b(n873) );
	nor2_1 U690 ( .x(n1083), .a(n4002), .b(___cell__39620_net143694) );
	nand2_2 U691 ( .x(n3665), .a(n1391), .b(n3451) );
	inv_5 U692 ( .x(n2022), .a(n1626) );
	inv_5 U693 ( .x(n3314), .a(n2136) );
	nand2_2 U694 ( .x(n3666), .a(n1256), .b(n2133) );
	oai211_1 U695 ( .x(n2046), .a(n1082), .b(n1664), .c(n2047), .d(n2048) );
	nand2_2 U696 ( .x(n2047), .a(n2193), .b(n3676) );
	inv_2 U697 ( .x(n3676), .a(n1460) );
	nand2i_2 U698 ( .x(n3670), .a(n1565), .b(n3278) );
	nand2i_2 U699 ( .x(n3671), .a(n1559), .b(n3622) );
	nand2i_2 U70 ( .x(n3293), .a(n1657), .b(n873) );
	inv_2 U700 ( .x(n1078), .a(N1805) );
	nor2_1 U701 ( .x(n1076), .a(n1077), .b(n1078) );
	nand2i_2 U702 ( .x(n3673), .a(n4005), .b(n1136) );
	nand2i_2 U703 ( .x(n3675), .a(n1608), .b(n3538) );
	nor2i_2 U704 ( .x(n1071), .a(n1042), .b(n1072) );
	inv_5 U705 ( .x(___cell__39620_net144303), .a(___cell__39620_net144302) );
	nor2i_0 U706 ( .x(n1074), .a(n914), .b(___cell__39620_net143694) );
	nor2i_1 U707 ( .x(n1073), .a(n1074), .b(___cell__39620_net143658) );
	nor2i_0 U708 ( .x(n1075), .a(N1706), .b(___cell__39620_net143660) );
	oai211_1 U709 ( .x(n2396), .a(n505), .b(___cell__39620_net144257), .c(n2397),
		.d(n2398) );
	inv_5 U71 ( .x(n873), .a(n1622) );
	nand2_2 U710 ( .x(n2398), .a(n2193), .b(n3768) );
	inv_2 U711 ( .x(n3768), .a(n1475) );
	aoi22_1 U712 ( .x(n2304), .a(n1714), .b(n2305), .c(n1249), .d(n2306) );
	oai21_1 U713 ( .x(n2324), .a(n816), .b(n3731), .c(n2304) );
	oai22_5 U714 ( .x(n2303), .a(n1585), .b(n836), .c(n3462), .d(n4125) );
	oai21_2 U715 ( .x(n2456), .a(n1564), .b(n1093), .c(n3761) );
	nand2i_2 U716 ( .x(n2409), .a(n621), .b(n2456) );
	oai21_1 U717 ( .x(n2455), .a(n1564), .b(n695), .c(___cell__39620_net147350) );
	nand2i_2 U718 ( .x(n2406), .a(n1747), .b(n1064) );
	oai21_1 U719 ( .x(n2405), .a(n4002), .b(___cell__39620_net144605), .c(n2406) );
	nand2i_2 U72 ( .x(n3305), .a(___cell__39620_net144257), .b(n873) );
	inv_2 U720 ( .x(n717), .a(net149122) );
	inv_2 U722 ( .x(n3409), .a(n2287) );
	aoi22_1 U723 ( .x(n2372), .a(n1714), .b(n2286), .c(n1249), .d(n2373) );
	nand2i_2 U724 ( .x(n3766), .a(n1747), .b(n530) );
	inv_0 U725 ( .x(n1747), .a(reg_out_B[29]) );
	inv_2 U726 ( .x(net151497), .a(IR_opcode_field[3]) );
	inv_2 U727 ( .x(___cell__39620_net144309), .a(___cell__39620_net144307) );
	or2_1 U728 ( .x(n495), .a(IR_opcode_field[0]), .b(IR_opcode_field[3]) );
	nand2i_2 U729 ( .x(___cell__39620_net144307), .a(n495), .b(___cell__39620_net143655) );
	nand2i_2 U73 ( .x(n3371), .a(n1561), .b(n926) );
	nand2_0 U730 ( .x(n2376), .a(Imm[29]), .b(n539) );
	inv_5 U731 ( .x(n1290), .a(n2633) );
	inv_5 U732 ( .x(n3427), .a(n3726) );
	oai21_1 U733 ( .x(n3727), .a(n891), .b(n3427), .c(n4140) );
	inv_12 U734 ( .x(n662), .a(n1182) );
	nor2_0 U735 ( .x(n1181), .a(n4140), .b(n1182) );
	nor2i_1 U736 ( .x(n782), .a(Imm[31]), .b(___cell__39620_net143693) );
	inv_2 U737 ( .x(n3520), .a(n3721) );
	inv_4 U738 ( .x(n3594), .a(n890) );
	oai21_1 U739 ( .x(n2274), .a(n1648), .b(n1281), .c(n2275) );
	nand2i_2 U74 ( .x(n3370), .a(n1564), .b(n874) );
	nand2i_4 U740 ( .x(n2280), .a(n3486), .b(n3487) );
	oai211_3 U741 ( .x(n2279), .a(n3397), .b(___cell__39620_net144317), .c(n3398),
		.d(n3399) );
	aoi22_1 U742 ( .x(n2282), .a(n1971), .b(n2283), .c(n1177), .d(n2284) );
	nand2_2 U743 ( .x(n2287), .a(n3473), .b(n3474) );
	aoi222_1 U744 ( .x(n2285), .a(n1256), .b(n2286), .c(n1150), .d(n2287),
		.e(n2273), .f(n644) );
	nand3_1 U745 ( .x(n734), .a(n733), .b(n1520), .c(___cell__39620_net144355) );
	aoi21_1 U746 ( .x(n517), .a(n671), .b(n3726), .c(n626) );
	nor2_0 U747 ( .x(n795), .a(net151904), .b(net149167) );
	inv_8 U748 ( .x(___cell__39620_net143326), .a(___cell__39620_net147731) );
	nand2_0 U749 ( .x(___cell__39620_net147296), .a(n1658), .b(n1641) );
	nor2_0 U75 ( .x(n2002), .a(IR_function_field[2]), .b(IR_function_field[3]) );
	inv_2 U750 ( .x(n835), .a(n3740) );
	nand2i_2 U751 ( .x(n3728), .a(n1085), .b(n621) );
	nand3i_1 U752 ( .x(n2289), .a(n1636), .b(n3728), .c(___cell__39620_net145472) );
	nand2i_2 U753 ( .x(n3736), .a(N70), .b(n530) );
	inv_2 U754 ( .x(n3737), .a(n3736) );
	inv_5 U755 ( .x(___cell__39620_net144344), .a(___cell__39620_net144340) );
	or3i_1 U756 ( .x(___cell__39620_net144350), .a(___cell__39620_net144344),
		.b(n783), .c(___cell__39620_net143653) );
	nand2i_2 U757 ( .x(n770), .a(___cell__39620_net144350), .b(___cell__39620_net147732) );
	nand2_2 U758 ( .x(n2258), .a(reg_out_A[31]), .b(Imm[31]) );
	exnor2_1 U759 ( .x(n1469), .a(reg_out_A[31]), .b(Imm[31]) );
	oai21_1 U760 ( .x(n2291), .a(n1469), .b(n690), .c(n2292) );
	aoi21_1 U761 ( .x(n2272), .a(n2273), .b(n609), .c(n1149) );
	nand2i_2 U762 ( .x(n3732), .a(n1634), .b(n2305) );
	nand4_1 U763 ( .x(n3730), .a(n2269), .b(n3729), .c(n2267), .d(n3375) );
	oai211_1 U764 ( .x(n2290), .a(n3731), .b(n1451), .c(n3732), .d(n2272) );
	nand2i_2 U765 ( .x(n2294), .a(N70), .b(n1064) );
	inv_4 U766 ( .x(n3735), .a(n1154) );
	nand2_2 U767 ( .x(n1155), .a(n2263), .b(n2264) );
	nand4i_1 U768 ( .x(n1154), .a(n2259), .b(n3733), .c(n2261), .d(n3734) );
	aoi21_1 U769 ( .x(n1153), .a(net149120), .b(n1154), .c(n1155) );
	nand2i_2 U77 ( .x(n1960), .a(reg_out_B[28]), .b(n1959) );
	nand3i_1 U770 ( .x(n1662), .a(n2004), .b(n1590), .c(n2005) );
	nand2_2 U771 ( .x(n2005), .a(n2003), .b(n3593) );
	aoi22_1 U772 ( .x(n2006), .a(n1526), .b(n1534), .c(n1540), .d(n1530) );
	inv_5 U773 ( .x(n3506), .a(n3695) );
	inv_2 U774 ( .x(n1927), .a(N1931) );
	nand2i_2 U775 ( .x(n3194), .a(n1927), .b(n3999) );
	nand2i_2 U776 ( .x(n3193), .a(n1928), .b(n1987) );
	inv_2 U777 ( .x(n1928), .a(N1798) );
	nand2i_3 U778 ( .x(n3986), .a(___cell__39620_net144345), .b(n1165) );
	nand2i_4 U779 ( .x(n3245), .a(n3185), .b(n3986) );
	inv_5 U78 ( .x(n601), .a(reg_out_B[22]) );
	inv_2 U780 ( .x(n1926), .a(N1732) );
	nand2i_2 U781 ( .x(n3189), .a(n1926), .b(___cell__39620_net145150) );
	aoi21_1 U782 ( .x(n3188), .a(N1699), .b(___cell__39620_net145190), .c(n1420) );
	inv_2 U783 ( .x(n1925), .a(N1633) );
	oai211_1 U784 ( .x(n3187), .a(___cell__39620_net143872), .b(n1925), .c(n3188),
		.d(n3189) );
	nor2i_1 U785 ( .x(n3181), .a(n694), .b(n1657) );
	exnor2_1 U786 ( .x(n1517), .a(n917), .b(net149122) );
	inv_2 U787 ( .x(n3504), .a(n3279) );
	aoi22_1 U788 ( .x(n2808), .a(n1714), .b(n2809), .c(n1249), .d(n2130) );
	exnor2_1 U789 ( .x(n1518), .a(n816), .b(n917) );
	nand2i_2 U790 ( .x(n3432), .a(n1562), .b(n3622) );
	inv_2 U791 ( .x(n3557), .a(n3555) );
	nand2i_2 U792 ( .x(n3431), .a(n4003), .b(n3278) );
	oai221_1 U793 ( .x(n3177), .a(n3178), .b(n1687), .c(n1657), .d(n1093),
		.e(n3179) );
	nand2i_3 U794 ( .x(n3984), .a(n1451), .b(n3752) );
	nand2_2 U795 ( .x(n1660), .a(n701), .b(n1661) );
	nand2_0 U796 ( .x(n3218), .a(___cell__39620_net145617), .b(net149122) );
	nand2i_2 U797 ( .x(n3217), .a(n4019), .b(n3057) );
	nand2i_2 U798 ( .x(n1640), .a(net152465), .b(IR_opcode_field[1]) );
	aoi22_1 U799 ( .x(n3200), .a(n2079), .b(n3201), .c(n3202), .d(n917) );
	nand2i_2 U800 ( .x(n3201), .a(n622), .b(n3488) );
	inv_2 U801 ( .x(n3489), .a(n3201) );
	aoi22_1 U802 ( .x(n3199), .a(n2266), .b(n902), .c(n1066), .d(n2337) );
	inv_4 U803 ( .x(n3753), .a(n1738) );
	inv_2 U804 ( .x(n2335), .a(n1281) );
	inv_2 U805 ( .x(n599), .a(n696) );
	oai221_1 U806 ( .x(n3197), .a(n1417), .b(n1690), .c(n1657), .d(n1093),
		.e(n3198) );
	nand2i_2 U807 ( .x(n3985), .a(n1451), .b(n3755) );
	inv_2 U808 ( .x(n1543), .a(n1541) );
	nand2i_2 U809 ( .x(n1452), .a(n496), .b(n1543) );
	inv_8 U81 ( .x(n628), .a(n1561) );
	inv_2 U810 ( .x(n3612), .a(n3564) );
	inv_2 U811 ( .x(n3178), .a(n1966) );
	inv_2 U812 ( .x(n3344), .a(n3348) );
	or2_1 U813 ( .x(n522), .a(n569), .b(n1569) );
	inv_2 U814 ( .x(n3601), .a(n522) );
	inv_2 U815 ( .x(n3316), .a(n3320) );
	inv_2 U816 ( .x(n3326), .a(n3329) );
	inv_2 U817 ( .x(n3663), .a(n1458) );
	nand2_2 U818 ( .x(n2008), .a(n2193), .b(n3663) );
	aoi21_1 U819 ( .x(n1062), .a(n904), .b(n530), .c(n1064) );
	nand2_0 U82 ( .x(n3625), .a(___cell__39620_net144330), .b(reg_out_A[28]) );
	inv_2 U820 ( .x(n3621), .a(n3500) );
	inv_2 U821 ( .x(n3333), .a(n3338) );
	oai22_1 U822 ( .x(n3414), .a(n915), .b(n1649), .c(n508), .d(n815) );
	nand2i_2 U823 ( .x(n3586), .a(n1632), .b(n521) );
	nand2_1 U824 ( .x(n3587), .a(n1714), .b(n2187) );
	nand3_1 U825 ( .x(n2027), .a(n3587), .b(n3586), .c(n1998) );
	nand4_3 U826 ( .x(n3583), .a(n3582), .b(n3580), .c(n3579), .d(n3581) );
	nand2i_2 U827 ( .x(n3581), .a(n1625), .b(n3457) );
	ao22_5 U828 ( .x(n2233), .a(n3318), .b(n857), .c(n814), .d(n3584) );
	inv_5 U829 ( .x(n722), .a(n3317) );
	nand2_0 U83 ( .x(n3636), .a(___cell__39620_net144330), .b(reg_out_A[29]) );
	nand2i_2 U830 ( .x(n3590), .a(n1623), .b(n4127) );
	nand2i_2 U831 ( .x(n2031), .a(n4045), .b(n3057) );
	nand2i_2 U833 ( .x(n3659), .a(n1607), .b(n3655) );
	nand2i_2 U834 ( .x(n3660), .a(n4007), .b(n1349) );
	nand2i_2 U835 ( .x(n3661), .a(n1608), .b(n3658) );
	nor2i_3 U836 ( .x(n1048), .a(n1049), .b(n4005) );
	nand2i_2 U837 ( .x(n3650), .a(n4006), .b(n3475) );
	nor2i_3 U838 ( .x(n1046), .a(n1047), .b(n1043) );
	nand4i_2 U839 ( .x(n1054), .a(n1046), .b(n3651), .c(n3650), .d(n3649) );
	nor2i_1 U84 ( .x(n1280), .a(n583), .b(n1281) );
	nor2i_1 U840 ( .x(n1050), .a(n1051), .b(___cell__39620_net143658) );
	nor2i_1 U841 ( .x(n1052), .a(N1707), .b(___cell__39620_net143660) );
	inv_2 U842 ( .x(n3018), .a(n3956) );
	nand2i_2 U843 ( .x(n3956), .a(n703), .b(n3931) );
	nor2_1 U844 ( .x(n1347), .a(n679), .b(n4023) );
	nand4_1 U845 ( .x(n3056), .a(n3947), .b(n3946), .c(n3945), .d(n3944) );
	nand2i_2 U846 ( .x(n3017), .a(n784), .b(n3056) );
	nand2i_2 U847 ( .x(n3016), .a(n1658), .b(n3926) );
	inv_2 U848 ( .x(n713), .a(___cell__39620_net144062) );
	nand2i_4 U85 ( .x(n2128), .a(n547), .b(n3463) );
	aoi22_1 U850 ( .x(n2990), .a(___cell__39620_net144517), .b(n2991), .c(n1391),
		.d(n2992) );
	nand2i_2 U851 ( .x(n3943), .a(n1625), .b(n3069) );
	oai211_1 U852 ( .x(n3008), .a(n630), .b(___cell__39620_net144062), .c(n3943),
		.d(n2990) );
	nand2i_2 U853 ( .x(n3949), .a(n1634), .b(n3544) );
	nand2i_2 U854 ( .x(n3950), .a(n727), .b(n2851) );
	nand2i_2 U855 ( .x(n3951), .a(n1635), .b(n2852) );
	nand4_1 U856 ( .x(n3013), .a(n3951), .b(n3950), .c(n3949), .d(n3948) );
	aoi22_2 U857 ( .x(n2993), .a(n1714), .b(n2994), .c(n1256), .d(n2995) );
	nand2i_2 U858 ( .x(n3942), .a(n1632), .b(n3302) );
	inv_12 U859 ( .x(n3584), .a(n822) );
	aoi21_1 U86 ( .x(n2804), .a(n1289), .b(n2128), .c(n1280) );
	oai211_1 U860 ( .x(n3012), .a(n3355), .b(n1636), .c(n3942), .d(n2993) );
	inv_5 U861 ( .x(n3439), .a(n3606) );
	inv_2 U862 ( .x(n3955), .a(n1506) );
	nand2_2 U863 ( .x(n2997), .a(n2193), .b(n3955) );
	aoi21_1 U864 ( .x(n1346), .a(n609), .b(n530), .c(n1064) );
	oai211_1 U865 ( .x(n2996), .a(n1346), .b(n1874), .c(n2997), .d(n2998) );
	inv_0 U866 ( .x(n1358), .a(reg_out_B[14]) );
	inv_2 U867 ( .x(n1881), .a(N1845) );
	inv_2 U868 ( .x(n1341), .a(N1812) );
	nor2_1 U869 ( .x(n1340), .a(n1077), .b(n1341) );
	nand2i_2 U87 ( .x(n2340), .a(n1635), .b(n3196) );
	nand2i_2 U870 ( .x(n3952), .a(n1607), .b(n3790) );
	nand2i_3 U871 ( .x(n3954), .a(n1608), .b(n3648) );
	nand4i_1 U872 ( .x(n2988), .a(n1332), .b(n3954), .c(n3953), .d(n3952) );
	nor2i_1 U873 ( .x(n1336), .a(net151622), .b(n1585) );
	nor2i_1 U874 ( .x(n1335), .a(n1336), .b(___cell__39620_net143658) );
	nor2i_1 U875 ( .x(n1337), .a(N1713), .b(___cell__39620_net143660) );
	and4i_2 U876 ( .x(n766), .a(n568), .b(N3304), .c(___cell__39620_net144303),
		.d(n1619) );
	nor2_0 U877 ( .x(n1327), .a(n4002), .b(___cell__39620_net143962) );
	nand4_1 U878 ( .x(n3009), .a(n3917), .b(n3916), .c(n3915), .d(n3914) );
	nand4_1 U879 ( .x(n3931), .a(n3930), .b(n3929), .c(n3928), .d(n3927) );
	nand2i_2 U880 ( .x(n2974), .a(___cell__39620_net144406), .b(n3931) );
	nand4_1 U881 ( .x(n3926), .a(n3925), .b(n3924), .c(n3923), .d(n3922) );
	ao22_3 U882 ( .x(n2977), .a(n3903), .b(n700), .c(n3926), .d(n757) );
	nand2i_2 U883 ( .x(n2979), .a(n4001), .b(n3897) );
	nor2_1 U884 ( .x(n1328), .a(n679), .b(n4024) );
	oai211_1 U885 ( .x(n2958), .a(n1326), .b(n1866), .c(n2959), .d(n2960) );
	aoi21_1 U886 ( .x(n1326), .a(n893), .b(n530), .c(n1064) );
	nand2_2 U887 ( .x(n2959), .a(n2193), .b(n3941) );
	inv_2 U888 ( .x(n3941), .a(n1504) );
	nand2i_2 U889 ( .x(n3933), .a(n1565), .b(n3622) );
	inv_8 U89 ( .x(n939), .a(n938) );
	inv_2 U890 ( .x(n1870), .a(N1879) );
	nand2i_2 U891 ( .x(n2952), .a(n1870), .b(n3998) );
	aoi211_1 U892 ( .x(n2948), .a(N1648), .b(n809), .c(n1325), .d(___cell__39620_net146132) );
	nor2i_1 U893 ( .x(n1325), .a(N1714), .b(___cell__39620_net143660) );
	oai22_1 U894 ( .x(___cell__39620_net146132), .a(n783), .b(n734), .c(___cell__39620_net143658),
		.d(___cell__39620_net146131) );
	inv_2 U895 ( .x(n1869), .a(N1747) );
	nand2i_2 U896 ( .x(n2951), .a(n1869), .b(___cell__39620_net145150) );
	aoi22_1 U897 ( .x(n2953), .a(N1979), .b(___cell__39620_net145508), .c(N1846),
		.d(n4000) );
	nand2i_2 U898 ( .x(n2957), .a(n1872), .b(n1987) );
	inv_2 U899 ( .x(n1872), .a(N1813) );
	buf_2 U90 ( .x(net149106), .a(Imm[1]) );
	nand2i_2 U900 ( .x(n2955), .a(n1616), .b(n1339) );
	and3i_1 U901 ( .x(n2914), .a(n2913), .b(n2915), .c(n2916) );
	nand2i_2 U902 ( .x(n2916), .a(n1860), .b(___cell__39620_net145190) );
	inv_2 U903 ( .x(n1860), .a(N1715) );
	oai22_1 U904 ( .x(n2913), .a(___cell__39620_net143872), .b(n1859), .c(___cell__39620_net143658),
		.d(n2912) );
	inv_2 U905 ( .x(n1859), .a(N1649) );
	inv_2 U906 ( .x(n1862), .a(N1880) );
	nand2i_2 U907 ( .x(n2919), .a(n1862), .b(n944) );
	nor2i_1 U908 ( .x(n1316), .a(n694), .b(n734) );
	aoi22_1 U909 ( .x(n2924), .a(N1847), .b(n4000), .c(N1980), .d(___cell__39620_net145508) );
	nand2i_2 U91 ( .x(n3698), .a(n1644), .b(n530) );
	nand2i_2 U910 ( .x(n2923), .a(n1864), .b(n1987) );
	inv_2 U911 ( .x(n1864), .a(N1814) );
	nand2i_2 U912 ( .x(n2922), .a(n1166), .b(n1339) );
	nand2i_2 U913 ( .x(n2921), .a(n1616), .b(n1308) );
	aoi21_2 U914 ( .x(n2762), .a(n1177), .b(n2763), .c(n2630) );
	inv_2 U915 ( .x(n3618), .a(n3405) );
	oai211_3 U916 ( .x(n2902), .a(n3620), .b(n1565), .c(n3857), .d(n2762) );
	nand2i_2 U917 ( .x(n3865), .a(n1562), .b(n2629) );
	nand2i_2 U918 ( .x(n3866), .a(n1565), .b(n3606) );
	inv_1 U919 ( .x(n827), .a(n761) );
	inv_2 U92 ( .x(n911), .a(reg_out_A[5]) );
	nand2i_2 U920 ( .x(n2929), .a(n1064), .b(n3913) );
	nand2i_2 U921 ( .x(n2934), .a(n1626), .b(n3887) );
	nand2i_2 U922 ( .x(n2933), .a(n1566), .b(n3004) );
	inv_1 U923 ( .x(net156025), .a(net156024) );
	inv_2 U924 ( .x(n638), .a(net156025) );
	oai21_1 U925 ( .x(n2932), .a(n1501), .b(n690), .c(n2935) );
	nand2i_2 U926 ( .x(n3896), .a(n1623), .b(n3547) );
	inv_5 U927 ( .x(n2943), .a(n2911) );
	nand2i_2 U928 ( .x(n3876), .a(n719), .b(n2784) );
	oai22_1 U929 ( .x(n2945), .a(n1087), .b(n4025), .c(n1217), .d(n1417) );
	exnor2_1 U93 ( .x(n1512), .a(reg_out_B[12]), .b(n894) );
	nand2i_2 U930 ( .x(n3878), .a(n1636), .b(n2781) );
	ao21_2 U931 ( .x(n516), .a(n1267), .b(n2938), .c(n1320) );
	nor2_1 U932 ( .x(n1320), .a(___cell__39620_net143693), .b(___cell__39620_net143954) );
	nand2i_2 U933 ( .x(n3898), .a(n727), .b(n2994) );
	nand2i_2 U934 ( .x(n3899), .a(n1634), .b(n3302) );
	nand2i_2 U935 ( .x(n3900), .a(n1632), .b(n3381) );
	nand2i_2 U936 ( .x(n3850), .a(n4003), .b(n3059) );
	inv_2 U937 ( .x(n3609), .a(n3309) );
	nand2i_4 U938 ( .x(n3610), .a(n3609), .b(n3598) );
	inv_6 U939 ( .x(n2696), .a(n2864) );
	oai22_1 U94 ( .x(n2082), .a(n2083), .b(n1687), .c(n1584), .d(n1690) );
	aoi21_2 U940 ( .x(n2672), .a(n1177), .b(n2673), .c(n2630) );
	inv_2 U941 ( .x(n3597), .a(n3474) );
	oai211_3 U942 ( .x(n2864), .a(n3600), .b(n1565), .c(n3845), .d(n2672) );
	aoai211_1 U943 ( .x(n2743), .a(n1217), .b(n2744), .c(n1561), .d(n2740) );
	inv_2 U944 ( .x(n2741), .a(n1491) );
	inv_2 U945 ( .x(n2742), .a(n1492) );
	mux2_2 U946 ( .x(n2711), .d0(n3378), .sl(n816), .d1(n3382) );
	nand2i_2 U947 ( .x(n2755), .a(___cell__39620_net144765), .b(___cell__39620_net145617) );
	inv_2 U948 ( .x(n3527), .a(n3733) );
	nand2i_2 U949 ( .x(n3526), .a(n3527), .b(n3528) );
	exnor2_1 U95 ( .x(n1479), .a(n533), .b(n681) );
	oai22_1 U950 ( .x(n3379), .a(n1587), .b(n915), .c(n853), .d(n815) );
	aoi21_1 U951 ( .x(n2737), .a(n1714), .b(n2738), .c(n1248) );
	nand2i_2 U952 ( .x(n3852), .a(n1634), .b(n3550) );
	nand2_1 U953 ( .x(n3853), .a(n504), .b(n2477) );
	nand3_1 U954 ( .x(n3854), .a(n3853), .b(n3852), .c(n2737) );
	nand2i_2 U955 ( .x(n3851), .a(n1623), .b(n2854) );
	inv_5 U956 ( .x(n799), .a(Imm[3]) );
	nand2i_2 U957 ( .x(n3843), .a(n1623), .b(n2784) );
	nor2_1 U958 ( .x(n1254), .a(n1087), .b(n4028) );
	aoi22_1 U959 ( .x(n2689), .a(n2690), .b(n1249), .c(n504), .d(n2433) );
	exnor2_1 U96 ( .x(n1480), .a(n533), .b(reg_out_B[27]) );
	nand2i_2 U960 ( .x(n3844), .a(n1634), .b(n2781) );
	oai22_2 U961 ( .x(n2779), .a(n506), .b(n536), .c(n1586), .d(n1629) );
	aoi22_1 U962 ( .x(n2727), .a(n663), .b(Imm[5]), .c(n662), .d(n2600) );
	inv_2 U963 ( .x(n1819), .a(N1719) );
	nand2i_2 U964 ( .x(n2726), .a(n1819), .b(___cell__39620_net145190) );
	oai211_1 U965 ( .x(n3839), .a(n844), .b(n4005), .c(n2632), .d(n3838) );
	nand2i_2 U966 ( .x(n2725), .a(n1055), .b(n3839) );
	nor2i_1 U967 ( .x(n1253), .a(N1851), .b(n946) );
	oai211_3 U968 ( .x(n2733), .a(n3656), .b(n1043), .c(n3846), .d(n2675) );
	inv_2 U969 ( .x(n709), .a(n802) );
	inv_2 U97 ( .x(n1931), .a(N1863) );
	inv_4 U970 ( .x(n1822), .a(N1951) );
	inv_2 U971 ( .x(n2676), .a(n4006) );
	inv_0 U972 ( .x(n1843), .a(reg_out_B[19]) );
	inv_2 U973 ( .x(n605), .a(reg_out_B[19]) );
	inv_5 U974 ( .x(n3550), .a(n752) );
	nand2i_2 U975 ( .x(n3831), .a(n1632), .b(n3550) );
	inv_2 U976 ( .x(n3406), .a(n2284) );
	nand2_2 U977 ( .x(n3832), .a(n1714), .b(n2477) );
	nand2_2 U978 ( .x(n3833), .a(n1256), .b(n2738) );
	inv_2 U979 ( .x(n2565), .a(n2277) );
	nand2i_2 U98 ( .x(n3250), .a(n1931), .b(n3997) );
	inv_5 U980 ( .x(n3454), .a(n2280) );
	inv_2 U981 ( .x(n3565), .a(n3640) );
	nand2i_4 U982 ( .x(n3820), .a(n4010), .b(n2520) );
	inv_16 U984 ( .x(n836), .a(n3575) );
	inv_2 U985 ( .x(n3403), .a(n2779) );
	nand2_2 U986 ( .x(n3822), .a(n1256), .b(n2779) );
	nand2_2 U987 ( .x(n3823), .a(n504), .b(n2306) );
	nand2i_2 U988 ( .x(n3824), .a(n1632), .b(n2781) );
	inv_2 U989 ( .x(n3310), .a(n2271) );
	nand2_0 U99 ( .x(n1621), .a(net152465), .b(IR_opcode_field[1]) );
	inv_2 U990 ( .x(n3534), .a(n3533) );
	inv_2 U991 ( .x(n3380), .a(n3379) );
	inv_8 U992 ( .x(n1561), .a(reg_out_A[21]) );
	exnor2_1 U993 ( .x(n1488), .a(n636), .b(n829) );
	exnor2_1 U994 ( .x(n1487), .a(n636), .b(reg_out_B[23]) );
	inv_2 U995 ( .x(n620), .a(___cell__6067_net21981) );
	nand2i_2 U996 ( .x(n1536), .a(___cell__39620_net144175), .b(n1537) );
	nand2i_5 U997 ( .x(n685), .a(n3604), .b(n3598) );
	aoi21_1 U998 ( .x(n2628), .a(n1177), .b(n2629), .c(n2630) );
	nand2i_2 U999 ( .x(n3836), .a(n4004), .b(n2981) );
	EX_DW01_add_32_5_test_1 add_271 ( .A({ reg_out_A[31], reg_out_A[30], reg_out_A[29],
		reg_out_A[28], n537, reg_out_A[26], n590, reg_out_A[24], n634, n686,
		reg_out_A[21], n749, reg_out_A[19], reg_out_A[18], reg_out_A[17], reg_out_A[16],
		n4016, n934, n930, reg_out_A[12], reg_out_A[11], reg_out_A[10], reg_out_A[9],
		reg_out_A[8], reg_out_A[7], n922, reg_out_A[5], reg_out_A[4], reg_out_A[3],
		n940, n832, n942}), .B({ Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26],
		n689, Imm[24], n829, n745, Imm[21], Imm[20], n684, Imm[18], Imm[17],
		Imm[16], Imm[15], Imm[14], Imm[13], n682, n753, Imm[10], Imm[9], Imm[8],
		Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], Imm[2], net149122, Imm[0]}),
		.CI(1'b0), .SUM({ N1729, N1728, N1727, N1726, N1725, N1724, N1723, N1722,
		N1721, N1720, N1719, N1718, N1717, N1716, N1715, N1714, N1713, N1712,
		N1711, N1710, N1709, N1708, N1707, N1706, N1705, N1704, N1703, N1702,
		N1701, N1700, N1699, N1698}), .CO() );
	EX_DW01_add_32_6_test_1 add_277 ( .A({ reg_out_A[31], reg_out_A[30], n539,
		reg_out_A[28], n533, reg_out_A[26], n590, reg_out_A[24], n634, n583,
		reg_out_A[21], n749, reg_out_A[19], reg_out_A[18], reg_out_A[17], reg_out_A[16],
		n4014, n934, n930, reg_out_A[12], reg_out_A[11], reg_out_A[10], reg_out_A[9],
		reg_out_A[8], reg_out_A[7], n921, reg_out_A[5], reg_out_A[4], reg_out_A[3],
		n939, n832, n943}), .B({ Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26],
		n689, Imm[24], n831, n745, Imm[21], Imm[20], Imm[19], Imm[18], Imm[17],
		Imm[16], Imm[15], Imm[14], Imm[13], Imm[12], Imm[11], Imm[10], Imm[9],
		Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], Imm[2], net149121, Imm[0]}),
		.CI(1'b0), .SUM({ N1762, N1761, N1760, N1759, N1758, N1757, N1756, N1755,
		N1754, N1753, N1752, N1751, N1750, N1749, N1748, N1747, N1746, N1745,
		N1744, N1743, N1742, N1741, N1740, N1739, N1738, N1737, N1736, N1735,
		N1734, N1733, N1732, N1731}), .CO() );
	EX_DW01_add_32_4_test_1 add_289 ( .A({ reg_out_A[31], reg_out_A[30], reg_out_A[29],
		reg_out_A[28], n537, reg_out_A[26], n590, reg_out_A[24], n636, n583,
		reg_out_A[21], reg_out_A[20], reg_out_A[19], reg_out_A[18], reg_out_A[17],
		reg_out_A[16], n608, n934, n930, reg_out_A[12], reg_out_A[11], reg_out_A[10],
		reg_out_A[9], reg_out_A[8], reg_out_A[7], n922, reg_out_A[5], reg_out_A[4],
		reg_out_A[3], n940, n832, n943}), .B({ Imm[31], Imm[30], Imm[29], Imm[28],
		n681, Imm[26], n689, Imm[24], n831, n745, Imm[21], Imm[20], Imm[19],
		Imm[18], Imm[17], Imm[16], Imm[15], Imm[14], Imm[13], Imm[12], Imm[11],
		Imm[10], Imm[9], Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], Imm[2],
		net149121, Imm[0]}), .CI(1'b0), .SUM({ N1828, N1827, N1826, N1825, N1824,
		N1823, N1822, N1821, N1820, N1819, N1818, N1817, N1816, N1815, N1814,
		N1813, N1812, N1811, N1810, N1809, N1808, N1807, N1806, N1805, N1804,
		N1803, N1802, N1801, N1800, N1799, N1798, N1797}), .CO() );
	EX_DW01_add_32_3_test_1 add_295 ( .A({ reg_out_A[31], n535, n539, n538,
		n533, reg_out_A[26], n590, reg_out_A[24], n636, n687, reg_out_A[21],
		reg_out_A[20], reg_out_A[19], reg_out_A[18], n863, reg_out_A[16], n4014,
		n933, n930, reg_out_A[12], reg_out_A[11], reg_out_A[10], reg_out_A[9],
		reg_out_A[8], reg_out_A[7], n936, reg_out_A[5], reg_out_A[4], reg_out_A[3],
		n940, n603, n942}), .B({ Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26],
		n689, Imm[24], n831, n745, Imm[21], Imm[20], Imm[19], Imm[18], Imm[17],
		Imm[16], Imm[15], Imm[14], Imm[13], Imm[12], Imm[11], Imm[10], Imm[9],
		Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], Imm[2], net149106, Imm[0]}),
		.CI(1'b0), .SUM({ N1861, N1860, N1859, N1858, N1857, N1856, N1855, N1854,
		N1853, N1852, N1851, N1850, N1849, N1848, N1847, N1846, N1845, N1844,
		N1843, N1842, N1841, N1840, N1839, N1838, N1837, N1836, N1835, N1834,
		N1833, N1832, N1831, N1830}), .CO() );
	EX_DW01_add_32_7_test_1 add_301 ( .A({ reg_out_A[31], reg_out_A[30], n539,
		n538, n533, n540, n590, reg_out_A[24], n636, n686, reg_out_A[21], n749,
		reg_out_A[19], reg_out_A[18], reg_out_A[17], reg_out_A[16], n602, n933,
		n930, reg_out_A[12], reg_out_A[11], reg_out_A[10], reg_out_A[9], reg_out_A[8],
		reg_out_A[7], n838, reg_out_A[5], reg_out_A[4], reg_out_A[3], n692, n603,
		n942}), .B({ Imm[31], Imm[30], Imm[29], Imm[28], n681, Imm[26], n689,
		Imm[24], n829, n745, Imm[21], n551, Imm[19], Imm[18], Imm[17], Imm[16],
		Imm[15], Imm[14], Imm[13], Imm[12], Imm[11], Imm[10], Imm[9], Imm[8],
		Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], n637, net149120, Imm[0]}), .CI(1'b0),
		.SUM({ N1894, N1893, N1892, N1891, N1890, N1889, N1888, N1887, N1886,
		N1885, N1884, N1883, N1882, N1881, N1880, N1879, N1878, N1877, N1876,
		N1875, N1874, N1873, N1872, N1871, N1870, N1869, N1868, N1867, N1866,
		N1865, N1864, N1863}), .CO() );
	EX_DW01_add_32_1_test_1 add_310 ( .A({ reg_out_A[31], reg_out_A[30], reg_out_A[29],
		n538, n537, n540, n590, n541, n634, n686, n628, n749, n887, n910, n902,
		n893, n609, n934, n930, n894, reg_out_A[11], n908, n904, reg_out_A[8],
		reg_out_A[7], n921, n912, n834, n885, n940, n832, n943}), .B({ 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, net151622, net156363, n556, n682, n753, Imm[10], net149617,
		Imm[8], Imm[7], Imm[6], net151578, net151904, net149167, n637, net149122,
		Imm[0]}), .CI(1'b0), .SUM({ N1961, N1960, N1959, N1958, N1957, N1956,
		N1955, N1954, N1953, N1952, N1951, N1950, N1949, N1948, N1947, N1946,
		N1945, N1944, N1943, N1942, N1941, N1940, N1939, N1938, N1937, N1936,
		N1935, N1934, N1933, N1932, N1931, N1930}), .CO() );
	smlatnr_1 byte_reg__master ( .q(byte_reg__m2s), .qb(), .d(n4048), .sdi(ALU_result[31]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 byte_reg__slave ( .q(_byte), .qb(n4046), .d(byte_reg__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	EX_DW01_cmp2_32_3_test_1 gte_246 ( .A({ N70, reg_out_B[30], reg_out_B[29],
		reg_out_B[28], reg_out_B[27], reg_out_B[26], reg_out_B[25], reg_out_B[24],
		reg_out_B[23], reg_out_B[22], n566, reg_out_B[20], reg_out_B[19], reg_out_B[18],
		reg_out_B[17], reg_out_B[16], reg_out_B[15], reg_out_B[14], reg_out_B[13],
		reg_out_B[12], reg_out_B[11], reg_out_B[10], reg_out_B[9], reg_out_B[8],
		n4146, reg_out_B[6], reg_out_B[5], reg_out_B[4], reg_out_B[3], n815,
		n816, reg_out_B[0]}), .B({ N69, reg_out_A[30], reg_out_A[29], reg_out_A[28],
		n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634, n583, reg_out_A[21],
		n749, n887, n910, n902, n893, n4016, n644, n930, n894, n901, n908, n904,
		n914, n852, n838, n912, n834, reg_out_A[3], n692, n917, n942}), .LEQ(1'b1),
		.TC(1'b0), .LT_LE(N1407), .GE_GT() );
	EX_DW01_cmp2_32_0 gte_348 ( .A({ N144, Imm[30], Imm[29], Imm[28], n681,
		Imm[26], n689, Imm[24], n829, n745, Imm[21], n551, n684, n633, n640,
		n631, net151622, net156363, n556, n682, n753, Imm[10], net149617, net149628,
		Imm[7], n642, net151578, net151904, n527, n891, n694, net152465}), .B({
		N69, reg_out_A[30], reg_out_A[29], reg_out_A[28], n533, reg_out_A[26],
		n590, n541, n636, n583, reg_out_A[21], n749, n887, n910, n902, n893,
		n608, n644, n930, n894, n901, n908, n904, n914, n852, n838, n912, n834,
		n885, n692, n917, n942}), .LEQ(1'b1), .TC(1'b0), .LT_LE(N3029), .GE_GT() );
	EX_DW01_cmp2_32_5_test_1 lt_240 ( .A({ N69, reg_out_A[30], reg_out_A[29],
		reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634,
		n686, n628, n749, n887, n910, n902, n893, n609, n644, n919, n894, n901,
		n908, n904, n914, n852, n838, n912, n834, reg_out_A[3], n692, n917, n943}),
		.B({ N70, reg_out_B[30], reg_out_B[29], reg_out_B[28], reg_out_B[27],
		reg_out_B[26], reg_out_B[25], reg_out_B[24], reg_out_B[23], reg_out_B[22],
		n566, reg_out_B[20], reg_out_B[19], reg_out_B[18], reg_out_B[17], reg_out_B[16],
		reg_out_B[15], reg_out_B[14], reg_out_B[13], reg_out_B[12], reg_out_B[11],
		reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, reg_out_B[6], reg_out_B[5],
		reg_out_B[4], reg_out_B[3], n815, n816, reg_out_B[0]}), .LEQ(1'b0), .TC(1'b0),
		.LT_LE(N1392), .GE_GT() );
	EX_DW01_cmp2_32_2 lt_342 ( .A({ N69, reg_out_A[30], reg_out_A[29], reg_out_A[28],
		n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n635, n583, reg_out_A[21],
		n749, n887, n910, n902, n893, n602, n644, n919, n894, n901, n908, n904,
		n914, reg_out_A[7], n920, n912, n834, reg_out_A[3], n692, n917, n943}),
		.B({ N144, Imm[30], Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], n831,
		n745, Imm[21], n551, n684, n633, n640, n631, net151622, net156363, n629,
		n682, n753, n818, net149617, net149628, Imm[7], Imm[6], net151578, net151904,
		Imm[3], n891, net149120, net152465}), .LEQ(1'b0), .TC(1'b0), .LT_LE(N3014),
		.GE_GT() );
	EX_DW01_cmp2_32_4_test_1 lte_242 ( .A({ N69, reg_out_A[30], reg_out_A[29],
		reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n636,
		n686, reg_out_A[21], n749, n596, n910, n902, n893, n609, n644, n524,
		n894, n901, n908, n904, n914, n852, n922, n912, n834, reg_out_A[3], n692,
		n917, n943}), .B({ N70, reg_out_B[30], reg_out_B[29], reg_out_B[28],
		reg_out_B[27], reg_out_B[26], reg_out_B[25], reg_out_B[24], reg_out_B[23],
		reg_out_B[22], n566, reg_out_B[20], reg_out_B[19], reg_out_B[18], reg_out_B[17],
		reg_out_B[16], reg_out_B[15], reg_out_B[14], reg_out_B[13], reg_out_B[12],
		reg_out_B[11], reg_out_B[10], reg_out_B[9], reg_out_B[8], n4146, reg_out_B[6],
		reg_out_B[5], reg_out_B[4], reg_out_B[3], n815, n816, reg_out_B[0]}),
		.LEQ(1'b1), .TC(1'b0), .LT_LE(N1402), .GE_GT() );
	EX_DW01_cmp2_32_1 lte_344 ( .A({ N69, reg_out_A[30], reg_out_A[29], reg_out_A[28],
		n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634, n686, n628,
		n749, n887, n910, n902, n893, n609, n644, n524, n894, n901, n908, n904,
		n914, n852, n922, n912, n834, n885, n692, n917, n943}), .B({ N144, Imm[30],
		Imm[29], Imm[28], n681, Imm[26], n689, Imm[24], n829, n745, Imm[21],
		n551, n684, n633, n639, n631, net151622, Imm[14], Imm[13], Imm[12], n753,
		n818, net149617, net149628, Imm[7], n642, net151578, net151904, Imm[3],
		n891, net149120, net152465}), .LEQ(1'b1), .TC(1'b0), .LT_LE(N3024), .GE_GT() );
	smlatnr_1 mem_read_EX_reg__master ( .q(mem_read_EX_reg__m2s), .qb(), .d(n4202),
		.sdi(_byte), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 mem_read_EX_reg__slave ( .q(mem_read_EX), .qb(), .d(mem_read_EX_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 mem_to_reg_EX_reg__master ( .q(mem_to_reg_EX_reg__m2s), .qb(),
		.d(n4200), .sdi(mem_read_EX), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 mem_to_reg_EX_reg__slave ( .q(n4224), .qb(n4201), .d(mem_to_reg_EX_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 mem_write_EX_reg__master ( .q(mem_write_EX_reg__m2s), .qb(),
		.d(n4203), .sdi(n4201), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 mem_write_EX_reg__slave ( .q(mem_write_EX), .qb(), .d(mem_write_EX_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	EX_DW01_sub_32_2_test_1 r1860_0 ( .A({ reg_out_A[31], reg_out_A[30], n539,
		n538, n537, n540, n590, n541, n634, n583, n628, reg_out_A[20], reg_out_A[19],
		reg_out_A[18], n586, n893, n608, n934, n918, reg_out_A[12], reg_out_A[11],
		n908, reg_out_A[9], reg_out_A[8], reg_out_A[7], n838, reg_out_A[5], reg_out_A[4],
		reg_out_A[3], n939, n832, n943}), .B({ n4144, reg_out_B[30], reg_out_B[29],
		reg_out_B[28], reg_out_B[27], reg_out_B[26], reg_out_B[25], reg_out_B[24],
		reg_out_B[23], reg_out_B[22], n567, reg_out_B[20], reg_out_B[19], reg_out_B[18],
		reg_out_B[17], reg_out_B[16], reg_out_B[15], reg_out_B[14], reg_out_B[13],
		reg_out_B[12], reg_out_B[11], reg_out_B[10], reg_out_B[9], reg_out_B[8],
		n4146, reg_out_B[6], reg_out_B[5], reg_out_B[4], reg_out_B[3], reg_out_B[2],
		reg_out_B[1], reg_out_B[0]}), .CI(1'b0), .DIFF({ N371, N370, N369, N368,
		N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, N356,
		N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, N344,
		N343, N342, N341, N340}), .CO() );
	EX_DW01_add_32_2_test_1 r1865_0 ( .A({ reg_out_A[31], reg_out_A[30], n539,
		reg_out_A[28], reg_out_A[27], reg_out_A[26], reg_out_A[25], reg_out_A[24],
		n634, n687, reg_out_A[21], n749, reg_out_A[19], reg_out_A[18], reg_out_A[17],
		reg_out_A[16], n4016, n934, n918, reg_out_A[12], reg_out_A[11], reg_out_A[10],
		reg_out_A[9], reg_out_A[8], reg_out_A[7], n921, reg_out_A[5], reg_out_A[4],
		reg_out_A[3], n939, n832, n943}), .B({ Imm[31], Imm[30], Imm[29], Imm[28],
		n681, Imm[26], n689, Imm[24], n829, n745, Imm[21], n551, Imm[19], Imm[18],
		Imm[17], Imm[16], Imm[15], Imm[14], Imm[13], Imm[12], Imm[11], Imm[10],
		Imm[9], Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], Imm[2], net149106,
		Imm[0]}), .CI(1'b0), .SUM({ N1663, N1662, N1661, N1660, N1659, N1658,
		N1657, N1656, N1655, N1654, N1653, N1652, N1651, N1650, N1649, N1648,
		N1647, N1646, N1645, N1644, N1643, N1642, N1641, N1640, N1639, N1638,
		N1637, N1636, N1635, N1634, N1633, N1632}), .CO() );
	EX_DW01_add_32_0_test_1 r247_0 ( .A({ reg_out_A[31], n535, reg_out_A[29],
		reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n634,
		n583, reg_out_A[21], reg_out_A[20], reg_out_A[19], reg_out_A[18], reg_out_A[17],
		reg_out_A[16], n608, n644, n930, n894, n901, n908, n904, n914, reg_out_A[7],
		n922, reg_out_A[5], reg_out_A[4], reg_out_A[3], n940, n832, n942}), .B({
		n4144, reg_out_B[30], reg_out_B[29], reg_out_B[28], reg_out_B[27], reg_out_B[26],
		reg_out_B[25], reg_out_B[24], reg_out_B[23], reg_out_B[22], n567, reg_out_B[20],
		reg_out_B[19], reg_out_B[18], reg_out_B[17], reg_out_B[16], reg_out_B[15],
		reg_out_B[14], reg_out_B[13], reg_out_B[12], reg_out_B[11], reg_out_B[10],
		reg_out_B[9], reg_out_B[8], n4146, reg_out_B[6], reg_out_B[5], reg_out_B[4],
		reg_out_B[3], reg_out_B[2], reg_out_B[1], reg_out_B[0]}), .CI(1'b0),
		.SUM({ N338, N337, N336, N335, N334, N333, N332, N331, N330, N329, N328,
		N327, N326, N325, N324, N323, N322, N321, N320, N319, N318, N317, N316,
		N315, N314, N313, N312, N311, N310, N309, N308, N307}), .CO() );
	smlatnr_1 reg_out_B_EX_reg_0__master ( .q(reg_out_B_EX_reg_0__m2s), .qb(),
		.d(n4212), .sdi(mem_write_EX), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_0__slave ( .q(reg_out_B_EX[0]), .qb(n4213), .d(reg_out_B_EX_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_10__master ( .q(reg_out_B_EX_reg_10__m2s), .qb(),
		.d(n4182), .sdi(n4209), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_10__slave ( .q(reg_out_B_EX[10]), .qb(n4183),
		.d(reg_out_B_EX_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_11__master ( .q(reg_out_B_EX_reg_11__m2s), .qb(),
		.d(n4214), .sdi(n4183), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_11__slave ( .q(reg_out_B_EX[11]), .qb(n4215),
		.d(reg_out_B_EX_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_12__master ( .q(reg_out_B_EX_reg_12__m2s), .qb(),
		.d(n4180), .sdi(n4215), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_12__slave ( .q(reg_out_B_EX[12]), .qb(n4181),
		.d(reg_out_B_EX_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_13__master ( .q(reg_out_B_EX_reg_13__m2s), .qb(),
		.d(n4216), .sdi(n4181), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_13__slave ( .q(reg_out_B_EX[13]), .qb(n4217),
		.d(reg_out_B_EX_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_14__master ( .q(reg_out_B_EX_reg_14__m2s), .qb(),
		.d(n4178), .sdi(n4217), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_14__slave ( .q(reg_out_B_EX[14]), .qb(n4179),
		.d(reg_out_B_EX_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_15__master ( .q(reg_out_B_EX_reg_15__m2s), .qb(),
		.d(n4158), .sdi(n4179), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_15__slave ( .q(reg_out_B_EX[15]), .qb(n4159),
		.d(reg_out_B_EX_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_16__master ( .q(reg_out_B_EX_reg_16__m2s), .qb(),
		.d(n4176), .sdi(n4159), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_16__slave ( .q(reg_out_B_EX[16]), .qb(n4177),
		.d(reg_out_B_EX_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_17__master ( .q(reg_out_B_EX_reg_17__m2s), .qb(),
		.d(n4222), .sdi(n4177), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_17__slave ( .q(reg_out_B_EX[17]), .qb(n4223),
		.d(reg_out_B_EX_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_18__master ( .q(reg_out_B_EX_reg_18__m2s), .qb(),
		.d(n4210), .sdi(n4223), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_18__slave ( .q(reg_out_B_EX[18]), .qb(n4211),
		.d(reg_out_B_EX_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_19__master ( .q(reg_out_B_EX_reg_19__m2s), .qb(),
		.d(n4174), .sdi(n4211), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_19__slave ( .q(reg_out_B_EX[19]), .qb(n4175),
		.d(reg_out_B_EX_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_1__master ( .q(reg_out_B_EX_reg_1__m2s), .qb(),
		.d(n4160), .sdi(n4213), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_1__slave ( .q(reg_out_B_EX[1]), .qb(n4161), .d(reg_out_B_EX_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_20__master ( .q(reg_out_B_EX_reg_20__m2s), .qb(),
		.d(n4218), .sdi(n4175), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_20__slave ( .q(reg_out_B_EX[20]), .qb(n4219),
		.d(reg_out_B_EX_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_21__master ( .q(reg_out_B_EX_reg_21__m2s), .qb(),
		.d(n4162), .sdi(n4219), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_21__slave ( .q(reg_out_B_EX[21]), .qb(n4163),
		.d(reg_out_B_EX_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_22__master ( .q(reg_out_B_EX_reg_22__m2s), .qb(),
		.d(n4204), .sdi(n4163), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_22__slave ( .q(reg_out_B_EX[22]), .qb(n4205),
		.d(reg_out_B_EX_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_23__master ( .q(reg_out_B_EX_reg_23__m2s), .qb(),
		.d(n4172), .sdi(n4205), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_23__slave ( .q(reg_out_B_EX[23]), .qb(n4173),
		.d(reg_out_B_EX_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_24__master ( .q(reg_out_B_EX_reg_24__m2s), .qb(),
		.d(n4156), .sdi(n4173), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_24__slave ( .q(reg_out_B_EX[24]), .qb(n4157),
		.d(reg_out_B_EX_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_25__master ( .q(reg_out_B_EX_reg_25__m2s), .qb(),
		.d(n4170), .sdi(n4157), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_25__slave ( .q(reg_out_B_EX[25]), .qb(n4171),
		.d(reg_out_B_EX_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_26__master ( .q(reg_out_B_EX_reg_26__m2s), .qb(),
		.d(n4206), .sdi(n4171), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_26__slave ( .q(reg_out_B_EX[26]), .qb(n4207),
		.d(reg_out_B_EX_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_27__master ( .q(reg_out_B_EX_reg_27__m2s), .qb(),
		.d(n4168), .sdi(n4207), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_27__slave ( .q(reg_out_B_EX[27]), .qb(n4169),
		.d(reg_out_B_EX_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_28__master ( .q(reg_out_B_EX_reg_28__m2s), .qb(),
		.d(n4166), .sdi(n4169), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_28__slave ( .q(reg_out_B_EX[28]), .qb(n4167),
		.d(reg_out_B_EX_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_29__master ( .q(reg_out_B_EX_reg_29__m2s), .qb(),
		.d(n4220), .sdi(n4167), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_29__slave ( .q(reg_out_B_EX[29]), .qb(n4221),
		.d(reg_out_B_EX_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_2__master ( .q(reg_out_B_EX_reg_2__m2s), .qb(),
		.d(n4196), .sdi(n4161), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_2__slave ( .q(reg_out_B_EX[2]), .qb(n4197), .d(reg_out_B_EX_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_30__master ( .q(reg_out_B_EX_reg_30__m2s), .qb(),
		.d(n4164), .sdi(n4221), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_30__slave ( .q(reg_out_B_EX[30]), .qb(n4165),
		.d(reg_out_B_EX_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_31__master ( .q(reg_out_B_EX_reg_31__m2s), .qb(),
		.d(N3297), .sdi(n4165), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_EX_reg_31__slave ( .q(reg_out_B_EX[31]), .qb(n4150),
		.d(reg_out_B_EX_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_3__master ( .q(reg_out_B_EX_reg_3__m2s), .qb(),
		.d(n4194), .sdi(n4197), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_3__slave ( .q(reg_out_B_EX[3]), .qb(n4195), .d(reg_out_B_EX_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_4__master ( .q(reg_out_B_EX_reg_4__m2s), .qb(),
		.d(n4192), .sdi(n4195), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_4__slave ( .q(reg_out_B_EX[4]), .qb(n4193), .d(reg_out_B_EX_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_5__master ( .q(reg_out_B_EX_reg_5__m2s), .qb(),
		.d(n4190), .sdi(n4193), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_5__slave ( .q(reg_out_B_EX[5]), .qb(n4191), .d(reg_out_B_EX_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_6__master ( .q(reg_out_B_EX_reg_6__m2s), .qb(),
		.d(n4188), .sdi(n4191), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_6__slave ( .q(reg_out_B_EX[6]), .qb(n4189), .d(reg_out_B_EX_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_7__master ( .q(reg_out_B_EX_reg_7__m2s), .qb(),
		.d(n4186), .sdi(n4189), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_7__slave ( .q(reg_out_B_EX[7]), .qb(n4187), .d(reg_out_B_EX_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_8__master ( .q(reg_out_B_EX_reg_8__m2s), .qb(),
		.d(n4184), .sdi(n4187), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_8__slave ( .q(reg_out_B_EX[8]), .qb(n4185), .d(reg_out_B_EX_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_EX_reg_9__master ( .q(reg_out_B_EX_reg_9__m2s), .qb(),
		.d(n4208), .sdi(n4185), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n543),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_EX_reg_9__slave ( .q(reg_out_B_EX[9]), .qb(n4209), .d(reg_out_B_EX_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n543), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_write_EX_reg__master ( .q(reg_write_EX_reg__m2s), .qb(),
		.d(n4198), .sdi(n4150), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4017),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_write_EX_reg__slave ( .q(reg_write_EX), .qb(n4199), .d(reg_write_EX_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4017), .glob_g(global_g2), .sync_sel(sync_sel) );
	EX_DW01_sub_32_0_test_1 sub_312 ( .A({ reg_out_A[31], reg_out_A[30], reg_out_A[29],
		reg_out_A[28], n533, reg_out_A[26], reg_out_A[25], reg_out_A[24], n636,
		n686, reg_out_A[21], reg_out_A[20], reg_out_A[19], reg_out_A[18], n902,
		n893, n602, n934, n930, reg_out_A[12], reg_out_A[11], reg_out_A[10],
		reg_out_A[9], reg_out_A[8], reg_out_A[7], n922, reg_out_A[5], reg_out_A[4],
		reg_out_A[3], n940, n917, n943}), .B({ Imm[31], Imm[30], Imm[29], Imm[28],
		n681, Imm[26], n689, Imm[24], n829, n745, Imm[21], Imm[20], n684, Imm[18],
		n640, n631, net151622, net156363, Imm[13], Imm[12], n753, Imm[10], Imm[9],
		Imm[8], Imm[7], Imm[6], Imm[5], Imm[4], Imm[3], n637, n694, net152465}),
		.CI(1'b0), .DIFF({ N1994, N1993, N1992, N1991, N1990, N1989, N1988, N1987,
		N1986, N1985, N1984, N1983, N1982, N1981, N1980, N1979, N1978, N1977,
		N1976, N1975, N1974, N1973, N1972, N1971, N1970, N1969, N1968, N1967,
		N1966, N1965, N1964, N1963}), .CO() );
	EX_DW01_sub_32_1_test_1 sub_314 ( .A({ reg_out_A[31], reg_out_A[30], reg_out_A[29],
		n538, n533, n540, n590, n541, n636, n583, n628, n749, n887, n910, n902,
		n893, n608, n934, n930, reg_out_A[12], n901, reg_out_A[10], n904, n914,
		reg_out_A[7], n921, n912, n834, n885, n692, n917, n943}), .B({ 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, net151622, net156363, Imm[13], Imm[12], n753, Imm[10],
		net149617, net149628, Imm[7], Imm[6], net151578, net151904, Imm[3], n637,
		net149120, net152465}), .CI(1'b0), .DIFF({ N2027, N2026, N2025, N2024,
		N2023, N2022, N2021, N2020, N2019, N2018, N2017, N2016, N2015, N2014,
		N2013, N2012, N2011, N2010, N2009, N2008, N2007, N2006, N2005, N2004,
		N2003, N2002, N2001, N2000, N1999, N1998, N1997, N1996}), .CO() );
	smlatnr_1 word_reg__master ( .q(word_reg__m2s), .qb(), .d(n4080), .sdi(n4199),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n542), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 word_reg__slave ( .q(word), .qb(n4047), .d(word_reg__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n542), .glob_g(global_g2), .sync_sel(sync_sel) );

endmodule


module DLX_sync_MUX_OP_32_5_32_2_test_1 (  D0_31, D0_30, D0_29, D0_28, D0_27,
	D0_26, D0_25, D0_24, D0_23, D0_22, D0_21, D0_20, D0_19, D0_18, D0_17,
	D0_16, D0_15, D0_14, D0_13, D0_12, D0_11, D0_10, D0_9, D0_8, D0_7, D0_6,
	D0_5, D0_4, D0_3, D0_2, D0_1, D0_0, D1_31, D1_30, D1_29, D1_28, D1_27,
	D1_26, D1_25, D1_24, D1_23, D1_22, D1_21, D1_20, D1_19, D1_18, D1_17,
	D1_16, D1_15, D1_14, D1_13, D1_12, D1_11, D1_10, D1_9, D1_8, D1_7, D1_6,
	D1_5, D1_4, D1_3, D1_2, D1_1, D1_0, D2_31, D2_30, D2_29, D2_28, D2_27,
	D2_26, D2_25, D2_24, D2_23, D2_22, D2_21, D2_20, D2_19, D2_18, D2_17,
	D2_16, D2_15, D2_14, D2_13, D2_12, D2_11, D2_10, D2_9, D2_8, D2_7, D2_6,
	D2_5, D2_4, D2_3, D2_2, D2_1, D2_0, D3_31, D3_30, D3_29, D3_28, D3_27,
	D3_26, D3_25, D3_24, D3_23, D3_22, D3_21, D3_20, D3_19, D3_18, D3_17,
	D3_16, D3_15, D3_14, D3_13, D3_12, D3_11, D3_10, D3_9, D3_8, D3_7, D3_6,
	D3_5, D3_4, D3_3, D3_2, D3_1, D3_0, D4_31, D4_30, D4_29, D4_28, D4_27,
	D4_26, D4_25, D4_24, D4_23, D4_22, D4_21, D4_20, D4_19, D4_18, D4_17,
	D4_16, D4_15, D4_14, D4_13, D4_12, D4_11, D4_10, D4_9, D4_8, D4_7, D4_6,
	D4_5, D4_4, D4_3, D4_2, D4_1, D4_0, D5_31, D5_30, D5_29, D5_28, D5_27,
	D5_26, D5_25, D5_24, D5_23, D5_22, D5_21, D5_20, D5_19, D5_18, D5_17,
	D5_16, D5_15, D5_14, D5_13, D5_12, D5_11, D5_10, D5_9, D5_8, D5_7, D5_6,
	D5_5, D5_4, D5_3, D5_2, D5_1, D5_0, D6_31, D6_30, D6_29, D6_28, D6_27,
	D6_26, D6_25, D6_24, D6_23, D6_22, D6_21, D6_20, D6_19, D6_18, D6_17,
	D6_16, D6_15, D6_14, D6_13, D6_12, D6_11, D6_10, D6_9, D6_8, D6_7, D6_6,
	D6_5, D6_4, D6_3, D6_2, D6_1, D6_0, D7_31, D7_30, D7_29, D7_28, D7_27,
	D7_26, D7_25, D7_24, D7_23, D7_22, D7_21, D7_20, D7_19, D7_18, D7_17,
	D7_16, D7_15, D7_14, D7_13, D7_12, D7_11, D7_10, D7_9, D7_8, D7_7, D7_6,
	D7_5, D7_4, D7_3, D7_2, D7_1, D7_0, D8_31, D8_30, D8_29, D8_28, D8_27,
	D8_26, D8_25, D8_24, D8_23, D8_22, D8_21, D8_20, D8_19, D8_18, D8_17,
	D8_16, D8_15, D8_14, D8_13, D8_12, D8_11, D8_10, D8_9, D8_8, D8_7, D8_6,
	D8_5, D8_4, D8_3, D8_2, D8_1, D8_0, D9_31, D9_30, D9_29, D9_28, D9_27,
	D9_26, D9_25, D9_24, D9_23, D9_22, D9_21, D9_20, D9_19, D9_18, D9_17,
	D9_16, D9_15, D9_14, D9_13, D9_12, D9_11, D9_10, D9_9, D9_8, D9_7, D9_6,
	D9_5, D9_4, D9_3, D9_2, D9_1, D9_0, D10_31, D10_30, D10_29, D10_28, D10_27,
	D10_26, D10_25, D10_24, D10_23, D10_22, D10_21, D10_20, D10_19, D10_18,
	D10_17, D10_16, D10_15, D10_14, D10_13, D10_12, D10_11, D10_10, D10_9,
	D10_8, D10_7, D10_6, D10_5, D10_4, D10_3, D10_2, D10_1, D10_0, D11_31,
	D11_30, D11_29, D11_28, D11_27, D11_26, D11_25, D11_24, D11_23, D11_22,
	D11_21, D11_20, D11_19, D11_18, D11_17, D11_16, D11_15, D11_14, D11_13,
	D11_12, D11_11, D11_10, D11_9, D11_8, D11_7, D11_6, D11_5, D11_4, D11_3,
	D11_2, D11_1, D11_0, D12_31, D12_30, D12_29, D12_28, D12_27, D12_26, D12_25,
	D12_24, D12_23, D12_22, D12_21, D12_20, D12_19, D12_18, D12_17, D12_16,
	D12_15, D12_14, D12_13, D12_12, D12_11, D12_10, D12_9, D12_8, D12_7, D12_6,
	D12_5, D12_4, D12_3, D12_2, D12_1, D12_0, D13_31, D13_30, D13_29, D13_28,
	D13_27, D13_26, D13_25, D13_24, D13_23, D13_22, D13_21, D13_20, D13_19,
	D13_18, D13_17, D13_16, D13_15, D13_14, D13_13, D13_12, D13_11, D13_10,
	D13_9, D13_8, D13_7, D13_6, D13_5, D13_4, D13_3, D13_2, D13_1, D13_0,
	D14_31, D14_30, D14_29, D14_28, D14_27, D14_26, D14_25, D14_24, D14_23,
	D14_22, D14_21, D14_20, D14_19, D14_18, D14_17, D14_16, D14_15, D14_14,
	D14_13, D14_12, D14_11, D14_10, D14_9, D14_8, D14_7, D14_6, D14_5, D14_4,
	D14_3, D14_2, D14_1, D14_0, D15_31, D15_30, D15_29, D15_28, D15_27, D15_26,
	D15_25, D15_24, D15_23, D15_22, D15_21, D15_20, D15_19, D15_18, D15_17,
	D15_16, D15_15, D15_14, D15_13, D15_12, D15_11, D15_10, D15_9, D15_8,
	D15_7, D15_6, D15_5, D15_4, D15_3, D15_2, D15_1, D15_0, D16_31, D16_30,
	D16_29, D16_28, D16_27, D16_26, D16_25, D16_24, D16_23, D16_22, D16_21,
	D16_20, D16_19, D16_18, D16_17, D16_16, D16_15, D16_14, D16_13, D16_12,
	D16_11, D16_10, D16_9, D16_8, D16_7, D16_6, D16_5, D16_4, D16_3, D16_2,
	D16_1, D16_0, D17_31, D17_30, D17_29, D17_28, D17_27, D17_26, D17_25,
	D17_24, D17_23, D17_22, D17_21, D17_20, D17_19, D17_18, D17_17, D17_16,
	D17_15, D17_14, D17_13, D17_12, D17_11, D17_10, D17_9, D17_8, D17_7, D17_6,
	D17_5, D17_4, D17_3, D17_2, D17_1, D17_0, D18_31, D18_30, D18_29, D18_28,
	D18_27, D18_26, D18_25, D18_24, D18_23, D18_22, D18_21, D18_20, D18_19,
	D18_18, D18_17, D18_16, D18_15, D18_14, D18_13, D18_12, D18_11, D18_10,
	D18_9, D18_8, D18_7, D18_6, D18_5, D18_4, D18_3, D18_2, D18_1, D18_0,
	D19_31, D19_30, D19_29, D19_28, D19_27, D19_26, D19_25, D19_24, D19_23,
	D19_22, D19_21, D19_20, D19_19, D19_18, D19_17, D19_16, D19_15, D19_14,
	D19_13, D19_12, D19_11, D19_10, D19_9, D19_8, D19_7, D19_6, D19_5, D19_4,
	D19_3, D19_2, D19_1, D19_0, D20_31, D20_30, D20_29, D20_28, D20_27, D20_26,
	D20_25, D20_24, D20_23, D20_22, D20_21, D20_20, D20_19, D20_18, D20_17,
	D20_16, D20_15, D20_14, D20_13, D20_12, D20_11, D20_10, D20_9, D20_8,
	D20_7, D20_6, D20_5, D20_4, D20_3, D20_2, D20_1, D20_0, D21_31, D21_30,
	D21_29, D21_28, D21_27, D21_26, D21_25, D21_24, D21_23, D21_22, D21_21,
	D21_20, D21_19, D21_18, D21_17, D21_16, D21_15, D21_14, D21_13, D21_12,
	D21_11, D21_10, D21_9, D21_8, D21_7, D21_6, D21_5, D21_4, D21_3, D21_2,
	D21_1, D21_0, D22_31, D22_30, D22_29, D22_28, D22_27, D22_26, D22_25,
	D22_24, D22_23, D22_22, D22_21, D22_20, D22_19, D22_18, D22_17, D22_16,
	D22_15, D22_14, D22_13, D22_12, D22_11, D22_10, D22_9, D22_8, D22_7, D22_6,
	D22_5, D22_4, D22_3, D22_2, D22_1, D22_0, D23_31, D23_30, D23_29, D23_28,
	D23_27, D23_26, D23_25, D23_24, D23_23, D23_22, D23_21, D23_20, D23_19,
	D23_18, D23_17, D23_16, D23_15, D23_14, D23_13, D23_12, D23_11, D23_10,
	D23_9, D23_8, D23_7, D23_6, D23_5, D23_4, D23_3, D23_2, D23_1, D23_0,
	D24_31, D24_30, D24_29, D24_28, D24_27, D24_26, D24_25, D24_24, D24_23,
	D24_22, D24_21, D24_20, D24_19, D24_18, D24_17, D24_16, D24_15, D24_14,
	D24_13, D24_12, D24_11, D24_10, D24_9, D24_8, D24_7, D24_6, D24_5, D24_4,
	D24_3, D24_2, D24_1, D24_0, D25_31, D25_30, D25_29, D25_28, D25_27, D25_26,
	D25_25, D25_24, D25_23, D25_22, D25_21, D25_20, D25_19, D25_18, D25_17,
	D25_16, D25_15, D25_14, D25_13, D25_12, D25_11, D25_10, D25_9, D25_8,
	D25_7, D25_6, D25_5, D25_4, D25_3, D25_2, D25_1, D25_0, D26_31, D26_30,
	D26_29, D26_28, D26_27, D26_26, D26_25, D26_24, D26_23, D26_22, D26_21,
	D26_20, D26_19, D26_18, D26_17, D26_16, D26_15, D26_14, D26_13, D26_12,
	D26_11, D26_10, D26_9, D26_8, D26_7, D26_6, D26_5, D26_4, D26_3, D26_2,
	D26_1, D26_0, D27_31, D27_30, D27_29, D27_28, D27_27, D27_26, D27_25,
	D27_24, D27_23, D27_22, D27_21, D27_20, D27_19, D27_18, D27_17, D27_16,
	D27_15, D27_14, D27_13, D27_12, D27_11, D27_10, D27_9, D27_8, D27_7, D27_6,
	D27_5, D27_4, D27_3, D27_2, D27_1, D27_0, D28_31, D28_30, D28_29, D28_28,
	D28_27, D28_26, D28_25, D28_24, D28_23, D28_22, D28_21, D28_20, D28_19,
	D28_18, D28_17, D28_16, D28_15, D28_14, D28_13, D28_12, D28_11, D28_10,
	D28_9, D28_8, D28_7, D28_6, D28_5, D28_4, D28_3, D28_2, D28_1, D28_0,
	D29_31, D29_30, D29_29, D29_28, D29_27, D29_26, D29_25, D29_24, D29_23,
	D29_22, D29_21, D29_20, D29_19, D29_18, D29_17, D29_16, D29_15, D29_14,
	D29_13, D29_12, D29_11, D29_10, D29_9, D29_8, D29_7, D29_6, D29_5, D29_4,
	D29_3, D29_2, D29_1, D29_0, D30_31, D30_30, D30_29, D30_28, D30_27, D30_26,
	D30_25, D30_24, D30_23, D30_22, D30_21, D30_20, D30_19, D30_18, D30_17,
	D30_16, D30_15, D30_14, D30_13, D30_12, D30_11, D30_10, D30_9, D30_8,
	D30_7, D30_6, D30_5, D30_4, D30_3, D30_2, D30_1, D30_0, D31_31, D31_30,
	D31_29, D31_28, D31_27, D31_26, D31_25, D31_24, D31_23, D31_22, D31_21,
	D31_20, D31_19, D31_18, D31_17, D31_16, D31_15, D31_14, D31_13, D31_12,
	D31_11, D31_10, D31_9, D31_8, D31_7, D31_6, D31_5, D31_4, D31_3, D31_2,
	D31_1, D31_0, S0, S1, S2, S3, S4, Z_31, Z_30, Z_29, Z_28, Z_27, Z_26,
	Z_25, Z_24, Z_23, Z_22, Z_21, Z_20, Z_19, Z_18, Z_17, Z_16, Z_15, Z_14,
	Z_13, Z_12, Z_11, Z_10, Z_9, Z_8, Z_7, Z_6, Z_5, Z_4, Z_3, Z_2, Z_1, Z_0 );

input  D0_31, D0_30, D0_29, D0_28, D0_27, D0_26, D0_25, D0_24, D0_23, D0_22,
	D0_21, D0_20, D0_19, D0_18, D0_17, D0_16, D0_15, D0_14, D0_13, D0_12,
	D0_11, D0_10, D0_9, D0_8, D0_7, D0_6, D0_5, D0_4, D0_3, D0_2, D0_1, D0_0,
	D1_31, D1_30, D1_29, D1_28, D1_27, D1_26, D1_25, D1_24, D1_23, D1_22,
	D1_21, D1_20, D1_19, D1_18, D1_17, D1_16, D1_15, D1_14, D1_13, D1_12,
	D1_11, D1_10, D1_9, D1_8, D1_7, D1_6, D1_5, D1_4, D1_3, D1_2, D1_1, D1_0,
	D2_31, D2_30, D2_29, D2_28, D2_27, D2_26, D2_25, D2_24, D2_23, D2_22,
	D2_21, D2_20, D2_19, D2_18, D2_17, D2_16, D2_15, D2_14, D2_13, D2_12,
	D2_11, D2_10, D2_9, D2_8, D2_7, D2_6, D2_5, D2_4, D2_3, D2_2, D2_1, D2_0,
	D3_31, D3_30, D3_29, D3_28, D3_27, D3_26, D3_25, D3_24, D3_23, D3_22,
	D3_21, D3_20, D3_19, D3_18, D3_17, D3_16, D3_15, D3_14, D3_13, D3_12,
	D3_11, D3_10, D3_9, D3_8, D3_7, D3_6, D3_5, D3_4, D3_3, D3_2, D3_1, D3_0,
	D4_31, D4_30, D4_29, D4_28, D4_27, D4_26, D4_25, D4_24, D4_23, D4_22,
	D4_21, D4_20, D4_19, D4_18, D4_17, D4_16, D4_15, D4_14, D4_13, D4_12,
	D4_11, D4_10, D4_9, D4_8, D4_7, D4_6, D4_5, D4_4, D4_3, D4_2, D4_1, D4_0,
	D5_31, D5_30, D5_29, D5_28, D5_27, D5_26, D5_25, D5_24, D5_23, D5_22,
	D5_21, D5_20, D5_19, D5_18, D5_17, D5_16, D5_15, D5_14, D5_13, D5_12,
	D5_11, D5_10, D5_9, D5_8, D5_7, D5_6, D5_5, D5_4, D5_3, D5_2, D5_1, D5_0,
	D6_31, D6_30, D6_29, D6_28, D6_27, D6_26, D6_25, D6_24, D6_23, D6_22,
	D6_21, D6_20, D6_19, D6_18, D6_17, D6_16, D6_15, D6_14, D6_13, D6_12,
	D6_11, D6_10, D6_9, D6_8, D6_7, D6_6, D6_5, D6_4, D6_3, D6_2, D6_1, D6_0,
	D7_31, D7_30, D7_29, D7_28, D7_27, D7_26, D7_25, D7_24, D7_23, D7_22,
	D7_21, D7_20, D7_19, D7_18, D7_17, D7_16, D7_15, D7_14, D7_13, D7_12,
	D7_11, D7_10, D7_9, D7_8, D7_7, D7_6, D7_5, D7_4, D7_3, D7_2, D7_1, D7_0,
	D8_31, D8_30, D8_29, D8_28, D8_27, D8_26, D8_25, D8_24, D8_23, D8_22,
	D8_21, D8_20, D8_19, D8_18, D8_17, D8_16, D8_15, D8_14, D8_13, D8_12,
	D8_11, D8_10, D8_9, D8_8, D8_7, D8_6, D8_5, D8_4, D8_3, D8_2, D8_1, D8_0,
	D9_31, D9_30, D9_29, D9_28, D9_27, D9_26, D9_25, D9_24, D9_23, D9_22,
	D9_21, D9_20, D9_19, D9_18, D9_17, D9_16, D9_15, D9_14, D9_13, D9_12,
	D9_11, D9_10, D9_9, D9_8, D9_7, D9_6, D9_5, D9_4, D9_3, D9_2, D9_1, D9_0,
	D10_31, D10_30, D10_29, D10_28, D10_27, D10_26, D10_25, D10_24, D10_23,
	D10_22, D10_21, D10_20, D10_19, D10_18, D10_17, D10_16, D10_15, D10_14,
	D10_13, D10_12, D10_11, D10_10, D10_9, D10_8, D10_7, D10_6, D10_5, D10_4,
	D10_3, D10_2, D10_1, D10_0, D11_31, D11_30, D11_29, D11_28, D11_27, D11_26,
	D11_25, D11_24, D11_23, D11_22, D11_21, D11_20, D11_19, D11_18, D11_17,
	D11_16, D11_15, D11_14, D11_13, D11_12, D11_11, D11_10, D11_9, D11_8,
	D11_7, D11_6, D11_5, D11_4, D11_3, D11_2, D11_1, D11_0, D12_31, D12_30,
	D12_29, D12_28, D12_27, D12_26, D12_25, D12_24, D12_23, D12_22, D12_21,
	D12_20, D12_19, D12_18, D12_17, D12_16, D12_15, D12_14, D12_13, D12_12,
	D12_11, D12_10, D12_9, D12_8, D12_7, D12_6, D12_5, D12_4, D12_3, D12_2,
	D12_1, D12_0, D13_31, D13_30, D13_29, D13_28, D13_27, D13_26, D13_25,
	D13_24, D13_23, D13_22, D13_21, D13_20, D13_19, D13_18, D13_17, D13_16,
	D13_15, D13_14, D13_13, D13_12, D13_11, D13_10, D13_9, D13_8, D13_7, D13_6,
	D13_5, D13_4, D13_3, D13_2, D13_1, D13_0, D14_31, D14_30, D14_29, D14_28,
	D14_27, D14_26, D14_25, D14_24, D14_23, D14_22, D14_21, D14_20, D14_19,
	D14_18, D14_17, D14_16, D14_15, D14_14, D14_13, D14_12, D14_11, D14_10,
	D14_9, D14_8, D14_7, D14_6, D14_5, D14_4, D14_3, D14_2, D14_1, D14_0,
	D15_31, D15_30, D15_29, D15_28, D15_27, D15_26, D15_25, D15_24, D15_23,
	D15_22, D15_21, D15_20, D15_19, D15_18, D15_17, D15_16, D15_15, D15_14,
	D15_13, D15_12, D15_11, D15_10, D15_9, D15_8, D15_7, D15_6, D15_5, D15_4,
	D15_3, D15_2, D15_1, D15_0, D16_31, D16_30, D16_29, D16_28, D16_27, D16_26,
	D16_25, D16_24, D16_23, D16_22, D16_21, D16_20, D16_19, D16_18, D16_17,
	D16_16, D16_15, D16_14, D16_13, D16_12, D16_11, D16_10, D16_9, D16_8,
	D16_7, D16_6, D16_5, D16_4, D16_3, D16_2, D16_1, D16_0, D17_31, D17_30,
	D17_29, D17_28, D17_27, D17_26, D17_25, D17_24, D17_23, D17_22, D17_21,
	D17_20, D17_19, D17_18, D17_17, D17_16, D17_15, D17_14, D17_13, D17_12,
	D17_11, D17_10, D17_9, D17_8, D17_7, D17_6, D17_5, D17_4, D17_3, D17_2,
	D17_1, D17_0, D18_31, D18_30, D18_29, D18_28, D18_27, D18_26, D18_25,
	D18_24, D18_23, D18_22, D18_21, D18_20, D18_19, D18_18, D18_17, D18_16,
	D18_15, D18_14, D18_13, D18_12, D18_11, D18_10, D18_9, D18_8, D18_7, D18_6,
	D18_5, D18_4, D18_3, D18_2, D18_1, D18_0, D19_31, D19_30, D19_29, D19_28,
	D19_27, D19_26, D19_25, D19_24, D19_23, D19_22, D19_21, D19_20, D19_19,
	D19_18, D19_17, D19_16, D19_15, D19_14, D19_13, D19_12, D19_11, D19_10,
	D19_9, D19_8, D19_7, D19_6, D19_5, D19_4, D19_3, D19_2, D19_1, D19_0,
	D20_31, D20_30, D20_29, D20_28, D20_27, D20_26, D20_25, D20_24, D20_23,
	D20_22, D20_21, D20_20, D20_19, D20_18, D20_17, D20_16, D20_15, D20_14,
	D20_13, D20_12, D20_11, D20_10, D20_9, D20_8, D20_7, D20_6, D20_5, D20_4,
	D20_3, D20_2, D20_1, D20_0, D21_31, D21_30, D21_29, D21_28, D21_27, D21_26,
	D21_25, D21_24, D21_23, D21_22, D21_21, D21_20, D21_19, D21_18, D21_17,
	D21_16, D21_15, D21_14, D21_13, D21_12, D21_11, D21_10, D21_9, D21_8,
	D21_7, D21_6, D21_5, D21_4, D21_3, D21_2, D21_1, D21_0, D22_31, D22_30,
	D22_29, D22_28, D22_27, D22_26, D22_25, D22_24, D22_23, D22_22, D22_21,
	D22_20, D22_19, D22_18, D22_17, D22_16, D22_15, D22_14, D22_13, D22_12,
	D22_11, D22_10, D22_9, D22_8, D22_7, D22_6, D22_5, D22_4, D22_3, D22_2,
	D22_1, D22_0, D23_31, D23_30, D23_29, D23_28, D23_27, D23_26, D23_25,
	D23_24, D23_23, D23_22, D23_21, D23_20, D23_19, D23_18, D23_17, D23_16,
	D23_15, D23_14, D23_13, D23_12, D23_11, D23_10, D23_9, D23_8, D23_7, D23_6,
	D23_5, D23_4, D23_3, D23_2, D23_1, D23_0, D24_31, D24_30, D24_29, D24_28,
	D24_27, D24_26, D24_25, D24_24, D24_23, D24_22, D24_21, D24_20, D24_19,
	D24_18, D24_17, D24_16, D24_15, D24_14, D24_13, D24_12, D24_11, D24_10,
	D24_9, D24_8, D24_7, D24_6, D24_5, D24_4, D24_3, D24_2, D24_1, D24_0,
	D25_31, D25_30, D25_29, D25_28, D25_27, D25_26, D25_25, D25_24, D25_23,
	D25_22, D25_21, D25_20, D25_19, D25_18, D25_17, D25_16, D25_15, D25_14,
	D25_13, D25_12, D25_11, D25_10, D25_9, D25_8, D25_7, D25_6, D25_5, D25_4,
	D25_3, D25_2, D25_1, D25_0, D26_31, D26_30, D26_29, D26_28, D26_27, D26_26,
	D26_25, D26_24, D26_23, D26_22, D26_21, D26_20, D26_19, D26_18, D26_17,
	D26_16, D26_15, D26_14, D26_13, D26_12, D26_11, D26_10, D26_9, D26_8,
	D26_7, D26_6, D26_5, D26_4, D26_3, D26_2, D26_1, D26_0, D27_31, D27_30,
	D27_29, D27_28, D27_27, D27_26, D27_25, D27_24, D27_23, D27_22, D27_21,
	D27_20, D27_19, D27_18, D27_17, D27_16, D27_15, D27_14, D27_13, D27_12,
	D27_11, D27_10, D27_9, D27_8, D27_7, D27_6, D27_5, D27_4, D27_3, D27_2,
	D27_1, D27_0, D28_31, D28_30, D28_29, D28_28, D28_27, D28_26, D28_25,
	D28_24, D28_23, D28_22, D28_21, D28_20, D28_19, D28_18, D28_17, D28_16,
	D28_15, D28_14, D28_13, D28_12, D28_11, D28_10, D28_9, D28_8, D28_7, D28_6,
	D28_5, D28_4, D28_3, D28_2, D28_1, D28_0, D29_31, D29_30, D29_29, D29_28,
	D29_27, D29_26, D29_25, D29_24, D29_23, D29_22, D29_21, D29_20, D29_19,
	D29_18, D29_17, D29_16, D29_15, D29_14, D29_13, D29_12, D29_11, D29_10,
	D29_9, D29_8, D29_7, D29_6, D29_5, D29_4, D29_3, D29_2, D29_1, D29_0,
	D30_31, D30_30, D30_29, D30_28, D30_27, D30_26, D30_25, D30_24, D30_23,
	D30_22, D30_21, D30_20, D30_19, D30_18, D30_17, D30_16, D30_15, D30_14,
	D30_13, D30_12, D30_11, D30_10, D30_9, D30_8, D30_7, D30_6, D30_5, D30_4,
	D30_3, D30_2, D30_1, D30_0, D31_31, D31_30, D31_29, D31_28, D31_27, D31_26,
	D31_25, D31_24, D31_23, D31_22, D31_21, D31_20, D31_19, D31_18, D31_17,
	D31_16, D31_15, D31_14, D31_13, D31_12, D31_11, D31_10, D31_9, D31_8,
	D31_7, D31_6, D31_5, D31_4, D31_3, D31_2, D31_1, D31_0, S0, S1, S2, S3,
	S4;
output  Z_31, Z_30, Z_29, Z_28, Z_27, Z_26, Z_25, Z_24, Z_23, Z_22, Z_21,
	Z_20, Z_19, Z_18, Z_17, Z_16, Z_15, Z_14, Z_13, Z_12, Z_11, Z_10, Z_9,
	Z_8, Z_7, Z_6, Z_5, Z_4, Z_3, Z_2, Z_1, Z_0;

wire n1, n10, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
	n11, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n12,
	n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n13, n130,
	n131, n132, n133, n134, n135, n136, n137, n138, n139, n14, n140, n141,
	n142, n143, n144, n145, n146, n147, n148, n149, n15, n150, n151, n152,
	n153, n154, n155, n156, n157, n158, n159, n16, n160, n161, n162, n163,
	n164, n165, n166, n167, n168, n169, n17, n170, n171, n172, n173, n174,
	n175, n176, n177, n178, n179, n18, n180, n181, n182, n183, n184, n185,
	n186, n187, n188, n189, n19, n190, n191, n192, n193, n194, n195, n196,
	n197, n198, n199, n2, n20, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n21, n210, n211, n212, n213, n214, n215, n216, n217, n218,
	n219, n22, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
	n23, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n24,
	n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n25, n250,
	n251, n252, n253, n254, n255, n256, n257, n258, n259, n26, n260, n261,
	n262, n263, n264, n265, n266, n267, n268, n269, n27, n270, n271, n272,
	n273, n274, n275, n276, n277, n278, n279, n28, n280, n281, n282, n283,
	n284, n285, n286, n287, n288, n289, n29, n290, n291, n292, n293, n294,
	n295, n296, n297, n298, n299, n3, n30, n300, n301, n302, n303, n304, n305,
	n306, n307, n308, n309, n31, n310, n311, n312, n313, n314, n315, n316,
	n317, n318, n319, n32, n320, n321, n322, n323, n324, n325, n326, n327,
	n328, n329, n33, n330, n331, n332, n333, n334, n335, n336, n337, n338,
	n339, n34, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
	n35, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n36,
	n360, n361, n362, n363, n364, n365, n366, n37, n38, n39, n4, n40, n41,
	n42, n43, n44, n45, n46, n47, n48, n49, n5, n50, n51, n52, n53, n54, n55,
	n56, n57, n58, n59, n6, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
	n7, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n8, n80, n81, n82,
	n83, n84, n85, n86, n87, n88, n89, n9, n90, n91, n92, n93, n94, n95, n96,
	n97, n98, n99;


	mux4_2 U1 ( .x(n111), .d0(D4_0), .d1(D12_0), .d2(D20_0), .d3(D28_0), .sl0(n11),
		.sl1(n32) );
	mux4_2 U10 ( .x(n250), .d0(D1_11), .d1(D9_11), .d2(D17_11), .d3(D25_11),
		.sl0(n11), .sl1(n38) );
	mux2_4 U100 ( .x(Z_20), .d0(n67), .sl(S0), .d1(n227) );
	mux2_4 U101 ( .x(Z_21), .d0(n68), .sl(S0), .d1(n228) );
	mux2_4 U102 ( .x(Z_22), .d0(n69), .sl(S0), .d1(n229) );
	mux2_4 U103 ( .x(Z_23), .d0(n70), .sl(S0), .d1(n230) );
	mux2_4 U104 ( .x(Z_24), .d0(n71), .sl(S0), .d1(n231) );
	mux2_4 U105 ( .x(Z_26), .d0(n73), .sl(S0), .d1(n233) );
	mux2_4 U106 ( .x(Z_28), .d0(n75), .sl(S0), .d1(n235) );
	mux2_4 U107 ( .x(Z_29), .d0(n76), .sl(S0), .d1(n236) );
	mux2_4 U108 ( .x(Z_30), .d0(n77), .sl(S0), .d1(n237) );
	mux2_4 U109 ( .x(Z_31), .d0(n78), .sl(S0), .d1(n238) );
	mux4_2 U11 ( .x(n122), .d0(D4_11), .d1(D12_11), .d2(D20_11), .d3(D28_11),
		.sl0(n24), .sl1(n32) );
	mux4_3 U110 ( .x(n47), .d0(n79), .d1(n143), .d2(n111), .d3(n175), .sl0(n4),
		.sl1(n1) );
	mux4_3 U111 ( .x(n48), .d0(n80), .d1(n144), .d2(n112), .d3(n176), .sl0(n10),
		.sl1(n1) );
	mux4_3 U112 ( .x(n49), .d0(n81), .d1(n145), .d2(n113), .d3(n177), .sl0(n4),
		.sl1(n2) );
	mux4_3 U113 ( .x(n50), .d0(n82), .d1(n146), .d2(n114), .d3(n178), .sl0(n4),
		.sl1(n2) );
	mux4_3 U114 ( .x(n52), .d0(n84), .d1(n148), .d2(n116), .d3(n180), .sl0(n4),
		.sl1(n2) );
	mux4_3 U115 ( .x(n53), .d0(n85), .d1(n149), .d2(n117), .d3(n181), .sl0(n4),
		.sl1(n2) );
	mux4_3 U116 ( .x(n54), .d0(n86), .d1(n150), .d2(n118), .d3(n182), .sl0(n3),
		.sl1(n2) );
	mux4_3 U117 ( .x(n55), .d0(n87), .d1(n151), .d2(n119), .d3(n183), .sl0(n3),
		.sl1(n1) );
	mux4_3 U118 ( .x(n56), .d0(n88), .d1(n152), .d2(n120), .d3(n184), .sl0(n4),
		.sl1(n2) );
	mux4_3 U119 ( .x(n57), .d0(n89), .d1(n153), .d2(n121), .d3(n185), .sl0(n4),
		.sl1(n1) );
	mux4_2 U12 ( .x(n154), .d0(D2_11), .d1(D10_11), .d2(D18_11), .d3(D26_11),
		.sl0(n15), .sl1(n34) );
	mux4_3 U120 ( .x(n58), .d0(n90), .d1(n154), .d2(n122), .d3(n186), .sl0(n3),
		.sl1(n1) );
	mux4_3 U121 ( .x(n60), .d0(n92), .d1(n156), .d2(n124), .d3(n188), .sl0(n3),
		.sl1(n2) );
	mux4_3 U122 ( .x(n61), .d0(n93), .d1(n157), .d2(n125), .d3(n189), .sl0(n9),
		.sl1(n2) );
	mux4_3 U123 ( .x(n62), .d0(n94), .d1(n158), .d2(n126), .d3(n190), .sl0(n4),
		.sl1(n2) );
	mux4_3 U124 ( .x(n63), .d0(n95), .d1(n159), .d2(n127), .d3(n191), .sl0(n9),
		.sl1(n2) );
	mux4_3 U125 ( .x(n64), .d0(n96), .d1(n160), .d2(n128), .d3(n192), .sl0(n4),
		.sl1(n2) );
	mux4_3 U126 ( .x(n66), .d0(n98), .d1(n162), .d2(n130), .d3(n194), .sl0(n9),
		.sl1(n1) );
	mux4_3 U127 ( .x(n67), .d0(n99), .d1(n163), .d2(n131), .d3(n195), .sl0(n3),
		.sl1(n2) );
	mux4_3 U128 ( .x(n68), .d0(n100), .d1(n164), .d2(n132), .d3(n196), .sl0(n3),
		.sl1(n1) );
	mux4_3 U129 ( .x(n69), .d0(n101), .d1(n165), .d2(n133), .d3(n197), .sl0(n9),
		.sl1(n1) );
	mux4_2 U13 ( .x(n90), .d0(D0_11), .d1(D8_11), .d2(D16_11), .d3(D24_11),
		.sl0(n23), .sl1(n30) );
	mux4_3 U130 ( .x(n71), .d0(n103), .d1(n167), .d2(n135), .d3(n199), .sl0(n4),
		.sl1(n1) );
	mux4_3 U131 ( .x(n72), .d0(n104), .d1(n168), .d2(n136), .d3(n200), .sl0(n9),
		.sl1(n2) );
	mux4_3 U132 ( .x(n73), .d0(n105), .d1(n169), .d2(n137), .d3(n201), .sl0(n10),
		.sl1(n1) );
	mux4_3 U133 ( .x(n75), .d0(n107), .d1(n171), .d2(n139), .d3(n203), .sl0(n10),
		.sl1(n1) );
	mux4_3 U134 ( .x(n76), .d0(n108), .d1(n172), .d2(n140), .d3(n204), .sl0(n10),
		.sl1(n1) );
	mux4_3 U135 ( .x(n78), .d0(n110), .d1(n174), .d2(n142), .d3(n206), .sl0(n9),
		.sl1(n1) );
	mux4_3 U136 ( .x(n80), .d0(D0_1), .d1(D8_1), .d2(D16_1), .d3(D24_1), .sl0(n11),
		.sl1(n30) );
	mux4_3 U137 ( .x(n81), .d0(D0_2), .d1(D8_2), .d2(D16_2), .d3(D24_2), .sl0(n26),
		.sl1(n30) );
	mux4_3 U138 ( .x(n82), .d0(D0_3), .d1(D8_3), .d2(D16_3), .d3(D24_3), .sl0(n26),
		.sl1(n30) );
	mux4_3 U139 ( .x(n83), .d0(D0_4), .d1(D8_4), .d2(D16_4), .d3(D24_4), .sl0(n17),
		.sl1(n30) );
	mux4_2 U14 ( .x(n136), .d0(D4_25), .d1(D12_25), .d2(D20_25), .d3(D28_25),
		.sl0(n15), .sl1(n33) );
	mux4_3 U140 ( .x(n84), .d0(D0_5), .d1(D8_5), .d2(D16_5), .d3(D24_5), .sl0(n19),
		.sl1(n30) );
	mux4_3 U141 ( .x(n85), .d0(D0_6), .d1(D8_6), .d2(D16_6), .d3(D24_6), .sl0(n23),
		.sl1(n30) );
	mux4_3 U142 ( .x(n86), .d0(D0_7), .d1(D8_7), .d2(D16_7), .d3(D24_7), .sl0(n17),
		.sl1(n30) );
	mux4_3 U143 ( .x(n88), .d0(D0_9), .d1(D8_9), .d2(D16_9), .d3(D24_9), .sl0(n18),
		.sl1(n30) );
	mux4_3 U144 ( .x(n89), .d0(D0_10), .d1(D8_10), .d2(D16_10), .d3(D24_10),
		.sl0(n28), .sl1(n30) );
	mux4_3 U145 ( .x(n92), .d0(D0_13), .d1(D8_13), .d2(D16_13), .d3(D24_13),
		.sl0(n17), .sl1(n30) );
	mux4_3 U146 ( .x(n93), .d0(D0_14), .d1(D8_14), .d2(D16_14), .d3(D24_14),
		.sl0(n23), .sl1(n30) );
	mux4_3 U147 ( .x(n94), .d0(D0_15), .d1(D8_15), .d2(D16_15), .d3(D24_15),
		.sl0(n29), .sl1(n30) );
	mux4_3 U148 ( .x(n95), .d0(D0_16), .d1(D8_16), .d2(D16_16), .d3(D24_16),
		.sl0(n11), .sl1(n31) );
	mux4_3 U149 ( .x(n96), .d0(D0_17), .d1(D8_17), .d2(D16_17), .d3(D24_17),
		.sl0(n20), .sl1(n31) );
	mux4_2 U15 ( .x(n168), .d0(D2_25), .d1(D10_25), .d2(D18_25), .d3(D26_25),
		.sl0(n19), .sl1(n35) );
	mux4_3 U150 ( .x(n97), .d0(D0_18), .d1(D8_18), .d2(D16_18), .d3(D24_18),
		.sl0(n17), .sl1(n31) );
	mux4_3 U151 ( .x(n98), .d0(D0_19), .d1(D8_19), .d2(D16_19), .d3(D24_19),
		.sl0(n18), .sl1(n31) );
	mux4_3 U152 ( .x(n99), .d0(D0_20), .d1(D8_20), .d2(D16_20), .d3(D24_20),
		.sl0(n23), .sl1(n31) );
	mux4_3 U153 ( .x(n100), .d0(D0_21), .d1(D8_21), .d2(D16_21), .d3(D24_21),
		.sl0(n18), .sl1(n31) );
	mux4_3 U154 ( .x(n101), .d0(D0_22), .d1(D8_22), .d2(D16_22), .d3(D24_22),
		.sl0(n23), .sl1(n31) );
	mux4_3 U155 ( .x(n102), .d0(D0_23), .d1(D8_23), .d2(D16_23), .d3(D24_23),
		.sl0(n28), .sl1(n31) );
	mux4_3 U156 ( .x(n103), .d0(D0_24), .d1(D8_24), .d2(D16_24), .d3(D24_24),
		.sl0(n16), .sl1(n31) );
	mux4_3 U157 ( .x(n104), .d0(D0_25), .d1(D8_25), .d2(D16_25), .d3(D24_25),
		.sl0(n29), .sl1(n31) );
	mux4_3 U158 ( .x(n105), .d0(D0_26), .d1(D8_26), .d2(D16_26), .d3(D24_26),
		.sl0(n23), .sl1(n31) );
	mux4_3 U159 ( .x(n106), .d0(D0_27), .d1(D8_27), .d2(D16_27), .d3(D24_27),
		.sl0(n23), .sl1(n31) );
	mux4_2 U16 ( .x(n123), .d0(D4_12), .d1(D12_12), .d2(D20_12), .d3(D28_12),
		.sl0(n15), .sl1(n32) );
	mux4_3 U160 ( .x(n107), .d0(D0_28), .d1(D8_28), .d2(D16_28), .d3(D24_28),
		.sl0(n23), .sl1(n31) );
	mux4_3 U161 ( .x(n108), .d0(D0_29), .d1(D8_29), .d2(D16_29), .d3(D24_29),
		.sl0(n18), .sl1(n31) );
	mux4_3 U162 ( .x(n109), .d0(D0_30), .d1(D8_30), .d2(D16_30), .d3(D24_30),
		.sl0(n23), .sl1(n31) );
	mux4_3 U163 ( .x(n110), .d0(D0_31), .d1(D8_31), .d2(D16_31), .d3(D24_31),
		.sl0(n23), .sl1(n31) );
	mux4_3 U164 ( .x(n112), .d0(D4_1), .d1(D12_1), .d2(D20_1), .d3(D28_1),
		.sl0(n16), .sl1(n32) );
	mux4_3 U165 ( .x(n113), .d0(D4_2), .d1(D12_2), .d2(D20_2), .d3(D28_2),
		.sl0(n19), .sl1(n32) );
	mux4_3 U166 ( .x(n114), .d0(D4_3), .d1(D12_3), .d2(D20_3), .d3(D28_3),
		.sl0(n23), .sl1(n32) );
	mux4_3 U167 ( .x(n115), .d0(D4_4), .d1(D12_4), .d2(D20_4), .d3(D28_4),
		.sl0(n19), .sl1(n32) );
	mux4_3 U168 ( .x(n116), .d0(D4_5), .d1(D12_5), .d2(D20_5), .d3(D28_5),
		.sl0(n11), .sl1(n32) );
	mux4_3 U169 ( .x(n117), .d0(D4_6), .d1(D12_6), .d2(D20_6), .d3(D28_6),
		.sl0(n19), .sl1(n32) );
	mux4_2 U17 ( .x(n91), .d0(D0_12), .d1(D8_12), .d2(D16_12), .d3(D24_12),
		.sl0(n17), .sl1(n30) );
	mux4_3 U170 ( .x(n118), .d0(D4_7), .d1(D12_7), .d2(D20_7), .d3(D28_7),
		.sl0(n29), .sl1(n32) );
	mux4_3 U171 ( .x(n120), .d0(D4_9), .d1(D12_9), .d2(D20_9), .d3(D28_9),
		.sl0(n11), .sl1(n32) );
	mux4_3 U172 ( .x(n121), .d0(D4_10), .d1(D12_10), .d2(D20_10), .d3(D28_10),
		.sl0(n24), .sl1(n32) );
	mux4_3 U173 ( .x(n124), .d0(D4_13), .d1(D12_13), .d2(D20_13), .d3(D28_13),
		.sl0(n26), .sl1(n32) );
	mux4_3 U174 ( .x(n125), .d0(D4_14), .d1(D12_14), .d2(D20_14), .d3(D28_14),
		.sl0(n15), .sl1(n32) );
	mux4_3 U175 ( .x(n126), .d0(D4_15), .d1(D12_15), .d2(D20_15), .d3(D28_15),
		.sl0(n24), .sl1(n32) );
	mux4_3 U176 ( .x(n127), .d0(D4_16), .d1(D12_16), .d2(D20_16), .d3(D28_16),
		.sl0(n24), .sl1(n33) );
	mux4_3 U177 ( .x(n128), .d0(D4_17), .d1(D12_17), .d2(D20_17), .d3(D28_17),
		.sl0(n15), .sl1(n33) );
	mux4_3 U178 ( .x(n129), .d0(D4_18), .d1(D12_18), .d2(D20_18), .d3(D28_18),
		.sl0(n24), .sl1(n33) );
	mux4_3 U179 ( .x(n130), .d0(D4_19), .d1(D12_19), .d2(D20_19), .d3(D28_19),
		.sl0(n29), .sl1(n33) );
	buf_8 U18 ( .x(n41), .a(S4) );
	mux4_3 U180 ( .x(n131), .d0(D4_20), .d1(D12_20), .d2(D20_20), .d3(D28_20),
		.sl0(n24), .sl1(n33) );
	mux4_3 U181 ( .x(n132), .d0(D4_21), .d1(D12_21), .d2(D20_21), .d3(D28_21),
		.sl0(n15), .sl1(n33) );
	mux4_3 U182 ( .x(n133), .d0(D4_22), .d1(D12_22), .d2(D20_22), .d3(D28_22),
		.sl0(n13), .sl1(n33) );
	mux4_3 U183 ( .x(n134), .d0(D4_23), .d1(D12_23), .d2(D20_23), .d3(D28_23),
		.sl0(n19), .sl1(n33) );
	mux4_3 U184 ( .x(n135), .d0(D4_24), .d1(D12_24), .d2(D20_24), .d3(D28_24),
		.sl0(n15), .sl1(n33) );
	mux4_3 U185 ( .x(n137), .d0(D4_26), .d1(D12_26), .d2(D20_26), .d3(D28_26),
		.sl0(n17), .sl1(n33) );
	mux4_3 U186 ( .x(n138), .d0(D4_27), .d1(D12_27), .d2(D20_27), .d3(D28_27),
		.sl0(n24), .sl1(n33) );
	mux4_3 U187 ( .x(n139), .d0(D4_28), .d1(D12_28), .d2(D20_28), .d3(D28_28),
		.sl0(n20), .sl1(n33) );
	mux4_3 U188 ( .x(n140), .d0(D4_29), .d1(D12_29), .d2(D20_29), .d3(D28_29),
		.sl0(n24), .sl1(n33) );
	mux4_3 U189 ( .x(n141), .d0(D4_30), .d1(D12_30), .d2(D20_30), .d3(D28_30),
		.sl0(n24), .sl1(n33) );
	buf_8 U19 ( .x(n35), .a(S4) );
	mux4_3 U190 ( .x(n142), .d0(D4_31), .d1(D12_31), .d2(D20_31), .d3(D28_31),
		.sl0(n15), .sl1(n33) );
	mux4_3 U191 ( .x(n144), .d0(D2_1), .d1(D10_1), .d2(D18_1), .d3(D26_1),
		.sl0(n26), .sl1(n34) );
	mux4_3 U192 ( .x(n145), .d0(D2_2), .d1(D10_2), .d2(D18_2), .d3(D26_2),
		.sl0(n24), .sl1(n34) );
	mux4_3 U193 ( .x(n146), .d0(D2_3), .d1(D10_3), .d2(D18_3), .d3(D26_3),
		.sl0(n24), .sl1(n34) );
	mux4_3 U194 ( .x(n147), .d0(D2_4), .d1(D10_4), .d2(D18_4), .d3(D26_4),
		.sl0(n15), .sl1(n34) );
	mux4_3 U195 ( .x(n148), .d0(D2_5), .d1(D10_5), .d2(D18_5), .d3(D26_5),
		.sl0(n24), .sl1(n34) );
	mux4_3 U196 ( .x(n149), .d0(D2_6), .d1(D10_6), .d2(D18_6), .d3(D26_6),
		.sl0(n24), .sl1(n34) );
	mux4_3 U197 ( .x(n150), .d0(D2_7), .d1(D10_7), .d2(D18_7), .d3(D26_7),
		.sl0(n20), .sl1(n34) );
	mux4_3 U198 ( .x(n151), .d0(D2_8), .d1(D10_8), .d2(D18_8), .d3(D26_8),
		.sl0(n25), .sl1(n34) );
	mux4_3 U199 ( .x(n152), .d0(D2_9), .d1(D10_9), .d2(D18_9), .d3(D26_9),
		.sl0(n15), .sl1(n34) );
	mux4_2 U2 ( .x(n143), .d0(D2_0), .d1(D10_0), .d2(D18_0), .d3(D26_0), .sl0(n15),
		.sl1(n34) );
	mux4_2 U20 ( .x(n211), .d0(n243), .d1(n307), .d2(n275), .d3(n339), .sl0(n4),
		.sl1(n2) );
	mux4_3 U200 ( .x(n153), .d0(D2_10), .d1(D10_10), .d2(D18_10), .d3(D26_10),
		.sl0(n20), .sl1(n34) );
	mux4_3 U201 ( .x(n155), .d0(D2_12), .d1(D10_12), .d2(D18_12), .d3(D26_12),
		.sl0(n25), .sl1(n34) );
	mux4_3 U202 ( .x(n156), .d0(D2_13), .d1(D10_13), .d2(D18_13), .d3(D26_13),
		.sl0(n13), .sl1(n34) );
	mux4_3 U203 ( .x(n157), .d0(D2_14), .d1(D10_14), .d2(D18_14), .d3(D26_14),
		.sl0(n20), .sl1(n34) );
	mux4_3 U204 ( .x(n158), .d0(D2_15), .d1(D10_15), .d2(D18_15), .d3(D26_15),
		.sl0(n28), .sl1(n34) );
	mux4_3 U205 ( .x(n159), .d0(D2_16), .d1(D10_16), .d2(D18_16), .d3(D26_16),
		.sl0(n15), .sl1(n35) );
	mux4_3 U206 ( .x(n160), .d0(D2_17), .d1(D10_17), .d2(D18_17), .d3(D26_17),
		.sl0(n25), .sl1(n35) );
	mux4_3 U207 ( .x(n161), .d0(D2_18), .d1(D10_18), .d2(D18_18), .d3(D26_18),
		.sl0(n13), .sl1(n35) );
	mux4_3 U208 ( .x(n162), .d0(D2_19), .d1(D10_19), .d2(D18_19), .d3(D26_19),
		.sl0(n25), .sl1(n35) );
	mux4_3 U209 ( .x(n163), .d0(D2_20), .d1(D10_20), .d2(D18_20), .d3(D26_20),
		.sl0(n25), .sl1(n35) );
	mux4_2 U21 ( .x(n51), .d0(n83), .d1(n147), .d2(n115), .d3(n179), .sl0(n3),
		.sl1(n2) );
	mux4_3 U210 ( .x(n164), .d0(D2_21), .d1(D10_21), .d2(D18_21), .d3(D26_21),
		.sl0(n15), .sl1(n35) );
	mux4_3 U211 ( .x(n165), .d0(D2_22), .d1(D10_22), .d2(D18_22), .d3(D26_22),
		.sl0(n15), .sl1(n35) );
	mux4_3 U212 ( .x(n166), .d0(D2_23), .d1(D10_23), .d2(D18_23), .d3(D26_23),
		.sl0(n18), .sl1(n35) );
	mux4_3 U213 ( .x(n167), .d0(D2_24), .d1(D10_24), .d2(D18_24), .d3(D26_24),
		.sl0(n25), .sl1(n35) );
	mux4_3 U214 ( .x(n169), .d0(D2_26), .d1(D10_26), .d2(D18_26), .d3(D26_26),
		.sl0(n25), .sl1(n35) );
	mux4_3 U215 ( .x(n170), .d0(D2_27), .d1(D10_27), .d2(D18_27), .d3(D26_27),
		.sl0(n20), .sl1(n35) );
	mux4_3 U216 ( .x(n171), .d0(D2_28), .d1(D10_28), .d2(D18_28), .d3(D26_28),
		.sl0(n14), .sl1(n35) );
	mux4_3 U217 ( .x(n172), .d0(D2_29), .d1(D10_29), .d2(D18_29), .d3(D26_29),
		.sl0(n14), .sl1(n35) );
	mux4_3 U218 ( .x(n173), .d0(D2_30), .d1(D10_30), .d2(D18_30), .d3(D26_30),
		.sl0(n14), .sl1(n35) );
	mux4_3 U219 ( .x(n174), .d0(D2_31), .d1(D10_31), .d2(D18_31), .d3(D26_31),
		.sl0(n25), .sl1(n35) );
	mux4_2 U22 ( .x(n214), .d0(n246), .d1(n310), .d2(n278), .d3(n342), .sl0(n3),
		.sl1(n2) );
	mux4_3 U220 ( .x(n175), .d0(D6_0), .d1(D14_0), .d2(D22_0), .d3(D30_0),
		.sl0(n25), .sl1(n36) );
	mux4_3 U221 ( .x(n176), .d0(D6_1), .d1(D14_1), .d2(D22_1), .d3(D30_1),
		.sl0(n29), .sl1(n36) );
	mux4_3 U222 ( .x(n177), .d0(D6_2), .d1(D14_2), .d2(D22_2), .d3(D30_2),
		.sl0(n25), .sl1(n36) );
	mux4_3 U223 ( .x(n178), .d0(D6_3), .d1(D14_3), .d2(D22_3), .d3(D30_3),
		.sl0(n25), .sl1(n36) );
	mux4_3 U224 ( .x(n179), .d0(D6_4), .d1(D14_4), .d2(D22_4), .d3(D30_4),
		.sl0(n14), .sl1(n36) );
	mux4_3 U225 ( .x(n180), .d0(D6_5), .d1(D14_5), .d2(D22_5), .d3(D30_5),
		.sl0(n29), .sl1(n36) );
	mux4_3 U226 ( .x(n181), .d0(D6_6), .d1(D14_6), .d2(D22_6), .d3(D30_6),
		.sl0(n14), .sl1(n36) );
	mux4_3 U227 ( .x(n182), .d0(D6_7), .d1(D14_7), .d2(D22_7), .d3(D30_7),
		.sl0(n14), .sl1(n36) );
	mux4_3 U228 ( .x(n184), .d0(D6_9), .d1(D14_9), .d2(D22_9), .d3(D30_9),
		.sl0(n18), .sl1(n36) );
	mux4_3 U229 ( .x(n185), .d0(D6_10), .d1(D14_10), .d2(D22_10), .d3(D30_10),
		.sl0(n19), .sl1(n36) );
	inv_3 U23 ( .x(Z_1), .a(n5) );
	mux4_3 U230 ( .x(n186), .d0(D6_11), .d1(D14_11), .d2(D22_11), .d3(D30_11),
		.sl0(n14), .sl1(n36) );
	mux4_3 U231 ( .x(n187), .d0(D6_12), .d1(D14_12), .d2(D22_12), .d3(D30_12),
		.sl0(n25), .sl1(n36) );
	mux4_3 U232 ( .x(n188), .d0(D6_13), .d1(D14_13), .d2(D22_13), .d3(D30_13),
		.sl0(n18), .sl1(n36) );
	mux4_3 U233 ( .x(n189), .d0(D6_14), .d1(D14_14), .d2(D22_14), .d3(D30_14),
		.sl0(n25), .sl1(n36) );
	mux4_3 U234 ( .x(n190), .d0(D6_15), .d1(D14_15), .d2(D22_15), .d3(D30_15),
		.sl0(n25), .sl1(n36) );
	mux4_3 U235 ( .x(n191), .d0(D6_16), .d1(D14_16), .d2(D22_16), .d3(D30_16),
		.sl0(n14), .sl1(n37) );
	mux4_3 U236 ( .x(n192), .d0(D6_17), .d1(D14_17), .d2(D22_17), .d3(D30_17),
		.sl0(n11), .sl1(n37) );
	mux4_3 U237 ( .x(n193), .d0(D6_18), .d1(D14_18), .d2(D22_18), .d3(D30_18),
		.sl0(n28), .sl1(n37) );
	mux4_3 U238 ( .x(n194), .d0(D6_19), .d1(D14_19), .d2(D22_19), .d3(D30_19),
		.sl0(n14), .sl1(n37) );
	mux4_3 U239 ( .x(n195), .d0(D6_20), .d1(D14_20), .d2(D22_20), .d3(D30_20),
		.sl0(n14), .sl1(n37) );
	mux4_3 U240 ( .x(n196), .d0(D6_21), .d1(D14_21), .d2(D22_21), .d3(D30_21),
		.sl0(n14), .sl1(n37) );
	mux4_3 U241 ( .x(n197), .d0(D6_22), .d1(D14_22), .d2(D22_22), .d3(D30_22),
		.sl0(n14), .sl1(n37) );
	mux4_3 U242 ( .x(n198), .d0(D6_23), .d1(D14_23), .d2(D22_23), .d3(D30_23),
		.sl0(n28), .sl1(n37) );
	mux4_3 U243 ( .x(n199), .d0(D6_24), .d1(D14_24), .d2(D22_24), .d3(D30_24),
		.sl0(n16), .sl1(n37) );
	mux4_3 U244 ( .x(n200), .d0(D6_25), .d1(D14_25), .d2(D22_25), .d3(D30_25),
		.sl0(n13), .sl1(n37) );
	mux4_3 U245 ( .x(n201), .d0(D6_26), .d1(D14_26), .d2(D22_26), .d3(D30_26),
		.sl0(n29), .sl1(n37) );
	mux4_3 U246 ( .x(n202), .d0(D6_27), .d1(D14_27), .d2(D22_27), .d3(D30_27),
		.sl0(n22), .sl1(n37) );
	mux4_3 U247 ( .x(n203), .d0(D6_28), .d1(D14_28), .d2(D22_28), .d3(D30_28),
		.sl0(n14), .sl1(n37) );
	mux4_3 U248 ( .x(n204), .d0(D6_29), .d1(D14_29), .d2(D22_29), .d3(D30_29),
		.sl0(n18), .sl1(n37) );
	mux4_3 U249 ( .x(n205), .d0(D6_30), .d1(D14_30), .d2(D22_30), .d3(D30_30),
		.sl0(n29), .sl1(n37) );
	mux4_2 U25 ( .x(n232), .d0(n264), .d1(n328), .d2(n296), .d3(n360), .sl0(n3),
		.sl1(n2) );
	mux4_3 U250 ( .x(n206), .d0(D6_31), .d1(D14_31), .d2(D22_31), .d3(D30_31),
		.sl0(n26), .sl1(n37) );
	mux4_3 U251 ( .x(n207), .d0(n239), .d1(n303), .d2(n271), .d3(n335), .sl0(n4),
		.sl1(n1) );
	mux4_3 U252 ( .x(n209), .d0(n241), .d1(n305), .d2(n273), .d3(n337), .sl0(n4),
		.sl1(n2) );
	mux4_3 U253 ( .x(n210), .d0(n242), .d1(n306), .d2(n274), .d3(n338), .sl0(n4),
		.sl1(n2) );
	mux4_3 U254 ( .x(n212), .d0(n244), .d1(n308), .d2(n276), .d3(n340), .sl0(n3),
		.sl1(n1) );
	mux4_3 U255 ( .x(n213), .d0(n245), .d1(n309), .d2(n277), .d3(n341), .sl0(n3),
		.sl1(n1) );
	mux4_3 U256 ( .x(n215), .d0(n247), .d1(n311), .d2(n279), .d3(n343), .sl0(n9),
		.sl1(n1) );
	mux4_3 U257 ( .x(n216), .d0(n248), .d1(n312), .d2(n280), .d3(n344), .sl0(n9),
		.sl1(n1) );
	mux4_3 U258 ( .x(n217), .d0(n249), .d1(n313), .d2(n281), .d3(n345), .sl0(n9),
		.sl1(n1) );
	mux4_3 U259 ( .x(n218), .d0(n250), .d1(n314), .d2(n282), .d3(n346), .sl0(n3),
		.sl1(n1) );
	mux4_2 U26 ( .x(n59), .d0(n91), .d1(n155), .d2(n123), .d3(n187), .sl0(n3),
		.sl1(n2) );
	mux4_3 U260 ( .x(n220), .d0(n252), .d1(n316), .d2(n284), .d3(n348), .sl0(n3),
		.sl1(n2) );
	mux4_3 U261 ( .x(n221), .d0(n253), .d1(n317), .d2(n285), .d3(n349), .sl0(n9),
		.sl1(n2) );
	mux4_3 U262 ( .x(n222), .d0(n254), .d1(n318), .d2(n286), .d3(n350), .sl0(n3),
		.sl1(n2) );
	mux4_3 U263 ( .x(n223), .d0(n255), .d1(n319), .d2(n287), .d3(n351), .sl0(n4),
		.sl1(n1) );
	mux4_3 U264 ( .x(n224), .d0(n256), .d1(n320), .d2(n288), .d3(n352), .sl0(n4),
		.sl1(n2) );
	mux4_3 U265 ( .x(n225), .d0(n257), .d1(n321), .d2(n289), .d3(n353), .sl0(n9),
		.sl1(n2) );
	mux4_3 U266 ( .x(n226), .d0(n258), .d1(n322), .d2(n290), .d3(n354), .sl0(n9),
		.sl1(n1) );
	mux4_3 U267 ( .x(n227), .d0(n259), .d1(n323), .d2(n291), .d3(n355), .sl0(n3),
		.sl1(n2) );
	mux4_3 U268 ( .x(n228), .d0(n260), .d1(n324), .d2(n292), .d3(n356), .sl0(n9),
		.sl1(n1) );
	mux4_3 U269 ( .x(n229), .d0(n261), .d1(n325), .d2(n293), .d3(n357), .sl0(n3),
		.sl1(n1) );
	mux4_2 U27 ( .x(n219), .d0(n251), .d1(n315), .d2(n283), .d3(n347), .sl0(n9),
		.sl1(n2) );
	mux4_3 U270 ( .x(n231), .d0(n263), .d1(n327), .d2(n295), .d3(n359), .sl0(n4),
		.sl1(n1) );
	mux4_3 U271 ( .x(n233), .d0(n265), .d1(n329), .d2(n297), .d3(n361), .sl0(n10),
		.sl1(n1) );
	mux4_3 U272 ( .x(n235), .d0(n267), .d1(n331), .d2(n299), .d3(n363), .sl0(n10),
		.sl1(n1) );
	mux4_3 U273 ( .x(n236), .d0(n268), .d1(n332), .d2(n300), .d3(n364), .sl0(n10),
		.sl1(n1) );
	mux4_3 U274 ( .x(n238), .d0(n270), .d1(n334), .d2(n302), .d3(n366), .sl0(n4),
		.sl1(n1) );
	mux4_3 U275 ( .x(n239), .d0(D1_0), .d1(D9_0), .d2(D17_0), .d3(D25_0), .sl0(n13),
		.sl1(n38) );
	mux4_3 U276 ( .x(n240), .d0(D1_1), .d1(D9_1), .d2(D17_1), .d3(D25_1), .sl0(n13),
		.sl1(n38) );
	mux4_3 U277 ( .x(n241), .d0(D1_2), .d1(D9_2), .d2(D17_2), .d3(D25_2), .sl0(n26),
		.sl1(n38) );
	mux4_3 U278 ( .x(n242), .d0(D1_3), .d1(D9_3), .d2(D17_3), .d3(D25_3), .sl0(n20),
		.sl1(n38) );
	mux4_3 U279 ( .x(n243), .d0(D1_4), .d1(D9_4), .d2(D17_4), .d3(D25_4), .sl0(n28),
		.sl1(n38) );
	mux2_2 U28 ( .x(Z_27), .d0(n74), .sl(S0), .d1(n234) );
	mux4_3 U280 ( .x(n244), .d0(D1_5), .d1(D9_5), .d2(D17_5), .d3(D25_5), .sl0(n29),
		.sl1(n38) );
	mux4_3 U281 ( .x(n245), .d0(D1_6), .d1(D9_6), .d2(D17_6), .d3(D25_6), .sl0(n28),
		.sl1(n38) );
	mux4_3 U282 ( .x(n246), .d0(D1_7), .d1(D9_7), .d2(D17_7), .d3(D25_7), .sl0(n26),
		.sl1(n38) );
	mux4_3 U283 ( .x(n247), .d0(D1_8), .d1(D9_8), .d2(D17_8), .d3(D25_8), .sl0(n29),
		.sl1(n38) );
	mux4_3 U284 ( .x(n248), .d0(D1_9), .d1(D9_9), .d2(D17_9), .d3(D25_9), .sl0(n17),
		.sl1(n38) );
	mux4_3 U285 ( .x(n249), .d0(D1_10), .d1(D9_10), .d2(D17_10), .d3(D25_10),
		.sl0(n19), .sl1(n38) );
	mux4_3 U286 ( .x(n251), .d0(D1_12), .d1(D9_12), .d2(D17_12), .d3(D25_12),
		.sl0(n20), .sl1(n38) );
	mux4_3 U287 ( .x(n252), .d0(D1_13), .d1(D9_13), .d2(D17_13), .d3(D25_13),
		.sl0(n26), .sl1(n38) );
	mux4_3 U288 ( .x(n253), .d0(D1_14), .d1(D9_14), .d2(D17_14), .d3(D25_14),
		.sl0(n29), .sl1(n38) );
	mux4_3 U289 ( .x(n254), .d0(D1_15), .d1(D9_15), .d2(D17_15), .d3(D25_15),
		.sl0(n20), .sl1(n38) );
	mux4_2 U29 ( .x(n74), .d0(n106), .d1(n170), .d2(n138), .d3(n202), .sl0(n9),
		.sl1(n2) );
	mux4_3 U290 ( .x(n255), .d0(D1_16), .d1(D9_16), .d2(D17_16), .d3(D25_16),
		.sl0(n26), .sl1(n39) );
	mux4_3 U291 ( .x(n256), .d0(D1_17), .d1(D9_17), .d2(D17_17), .d3(D25_17),
		.sl0(n29), .sl1(n39) );
	mux4_3 U292 ( .x(n257), .d0(D1_18), .d1(D9_18), .d2(D17_18), .d3(D25_18),
		.sl0(n19), .sl1(n39) );
	mux4_3 U293 ( .x(n258), .d0(D1_19), .d1(D9_19), .d2(D17_19), .d3(D25_19),
		.sl0(n16), .sl1(n39) );
	mux4_3 U294 ( .x(n259), .d0(D1_20), .d1(D9_20), .d2(D17_20), .d3(D25_20),
		.sl0(n17), .sl1(n39) );
	mux4_3 U295 ( .x(n260), .d0(D1_21), .d1(D9_21), .d2(D17_21), .d3(D25_21),
		.sl0(n28), .sl1(n39) );
	mux4_3 U296 ( .x(n261), .d0(D1_22), .d1(D9_22), .d2(D17_22), .d3(D25_22),
		.sl0(n19), .sl1(n39) );
	mux4_3 U297 ( .x(n262), .d0(D1_23), .d1(D9_23), .d2(D17_23), .d3(D25_23),
		.sl0(n13), .sl1(n39) );
	mux4_3 U298 ( .x(n263), .d0(D1_24), .d1(D9_24), .d2(D17_24), .d3(D25_24),
		.sl0(n26), .sl1(n39) );
	mux4_3 U299 ( .x(n264), .d0(D1_25), .d1(D9_25), .d2(D17_25), .d3(D25_25),
		.sl0(n25), .sl1(n39) );
	mux4_2 U3 ( .x(n79), .d0(D0_0), .d1(D8_0), .d2(D16_0), .d3(D24_0), .sl0(n17),
		.sl1(n30) );
	mux4_2 U30 ( .x(n234), .d0(n266), .d1(n330), .d2(n298), .d3(n362), .sl0(n4),
		.sl1(n2) );
	mux4_3 U300 ( .x(n265), .d0(D1_26), .d1(D9_26), .d2(D17_26), .d3(D25_26),
		.sl0(n13), .sl1(n39) );
	mux4_3 U301 ( .x(n266), .d0(D1_27), .d1(D9_27), .d2(D17_27), .d3(D25_27),
		.sl0(n16), .sl1(n39) );
	mux4_3 U302 ( .x(n267), .d0(D1_28), .d1(D9_28), .d2(D17_28), .d3(D25_28),
		.sl0(n20), .sl1(n39) );
	mux4_3 U303 ( .x(n268), .d0(D1_29), .d1(D9_29), .d2(D17_29), .d3(D25_29),
		.sl0(n13), .sl1(n39) );
	mux4_3 U304 ( .x(n269), .d0(D1_30), .d1(D9_30), .d2(D17_30), .d3(D25_30),
		.sl0(n21), .sl1(n39) );
	mux4_3 U305 ( .x(n270), .d0(D1_31), .d1(D9_31), .d2(D17_31), .d3(D25_31),
		.sl0(n19), .sl1(n39) );
	mux4_3 U306 ( .x(n271), .d0(D5_0), .d1(D13_0), .d2(D21_0), .d3(D29_0),
		.sl0(n20), .sl1(n40) );
	mux4_3 U307 ( .x(n272), .d0(D5_1), .d1(D13_1), .d2(D21_1), .d3(D29_1),
		.sl0(n11), .sl1(n40) );
	mux4_3 U308 ( .x(n273), .d0(D5_2), .d1(D13_2), .d2(D21_2), .d3(D29_2),
		.sl0(n13), .sl1(n40) );
	mux4_3 U309 ( .x(n274), .d0(D5_3), .d1(D13_3), .d2(D21_3), .d3(D29_3),
		.sl0(n11), .sl1(n40) );
	mux4_2 U31 ( .x(n65), .d0(n97), .d1(n161), .d2(n129), .d3(n193), .sl0(n3),
		.sl1(n2) );
	mux4_3 U310 ( .x(n275), .d0(D5_4), .d1(D13_4), .d2(D21_4), .d3(D29_4),
		.sl0(n21), .sl1(n40) );
	mux4_3 U311 ( .x(n276), .d0(D5_5), .d1(D13_5), .d2(D21_5), .d3(D29_5),
		.sl0(n18), .sl1(n40) );
	mux4_3 U312 ( .x(n277), .d0(D5_6), .d1(D13_6), .d2(D21_6), .d3(D29_6),
		.sl0(n17), .sl1(n40) );
	mux4_3 U313 ( .x(n278), .d0(D5_7), .d1(D13_7), .d2(D21_7), .d3(D29_7),
		.sl0(n21), .sl1(n40) );
	mux4_3 U314 ( .x(n280), .d0(D5_9), .d1(D13_9), .d2(D21_9), .d3(D29_9),
		.sl0(n12), .sl1(n40) );
	mux4_3 U315 ( .x(n281), .d0(D5_10), .d1(D13_10), .d2(D21_10), .d3(D29_10),
		.sl0(n12), .sl1(n40) );
	mux4_3 U316 ( .x(n283), .d0(D5_12), .d1(D13_12), .d2(D21_12), .d3(D29_12),
		.sl0(n21), .sl1(n40) );
	mux4_3 U317 ( .x(n284), .d0(D5_13), .d1(D13_13), .d2(D21_13), .d3(D29_13),
		.sl0(n21), .sl1(n40) );
	mux4_3 U318 ( .x(n285), .d0(D5_14), .d1(D13_14), .d2(D21_14), .d3(D29_14),
		.sl0(n27), .sl1(n40) );
	mux4_3 U319 ( .x(n286), .d0(D5_15), .d1(D13_15), .d2(D21_15), .d3(D29_15),
		.sl0(n12), .sl1(n40) );
	mux4_2 U32 ( .x(n230), .d0(n262), .d1(n326), .d2(n294), .d3(n358), .sl0(n3),
		.sl1(n2) );
	mux4_3 U320 ( .x(n287), .d0(D5_16), .d1(D13_16), .d2(D21_16), .d3(D29_16),
		.sl0(n12), .sl1(n41) );
	mux4_3 U321 ( .x(n288), .d0(D5_17), .d1(D13_17), .d2(D21_17), .d3(D29_17),
		.sl0(n21), .sl1(n41) );
	mux4_3 U322 ( .x(n289), .d0(D5_18), .d1(D13_18), .d2(D21_18), .d3(D29_18),
		.sl0(n12), .sl1(n41) );
	mux4_3 U323 ( .x(n290), .d0(D5_19), .d1(D13_19), .d2(D21_19), .d3(D29_19),
		.sl0(n27), .sl1(n41) );
	mux4_3 U324 ( .x(n291), .d0(D5_20), .d1(D13_20), .d2(D21_20), .d3(D29_20),
		.sl0(n21), .sl1(n41) );
	mux4_3 U325 ( .x(n292), .d0(D5_21), .d1(D13_21), .d2(D21_21), .d3(D29_21),
		.sl0(n27), .sl1(n41) );
	mux4_3 U326 ( .x(n293), .d0(D5_22), .d1(D13_22), .d2(D21_22), .d3(D29_22),
		.sl0(n27), .sl1(n41) );
	mux4_3 U327 ( .x(n294), .d0(D5_23), .d1(D13_23), .d2(D21_23), .d3(D29_23),
		.sl0(n12), .sl1(n41) );
	mux4_3 U328 ( .x(n295), .d0(D5_24), .d1(D13_24), .d2(D21_24), .d3(D29_24),
		.sl0(n27), .sl1(n41) );
	mux4_3 U329 ( .x(n296), .d0(D5_25), .d1(D13_25), .d2(D21_25), .d3(D29_25),
		.sl0(n27), .sl1(n41) );
	mux4_2 U33 ( .x(n70), .d0(n102), .d1(n166), .d2(n134), .d3(n198), .sl0(n3),
		.sl1(n2) );
	mux4_3 U330 ( .x(n297), .d0(D5_26), .d1(D13_26), .d2(D21_26), .d3(D29_26),
		.sl0(n27), .sl1(n41) );
	mux4_3 U331 ( .x(n298), .d0(D5_27), .d1(D13_27), .d2(D21_27), .d3(D29_27),
		.sl0(n27), .sl1(n41) );
	mux4_3 U332 ( .x(n299), .d0(D5_28), .d1(D13_28), .d2(D21_28), .d3(D29_28),
		.sl0(n27), .sl1(n41) );
	mux4_3 U333 ( .x(n300), .d0(D5_29), .d1(D13_29), .d2(D21_29), .d3(D29_29),
		.sl0(n21), .sl1(n41) );
	mux4_3 U334 ( .x(n301), .d0(D5_30), .d1(D13_30), .d2(D21_30), .d3(D29_30),
		.sl0(n21), .sl1(n41) );
	mux4_3 U335 ( .x(n302), .d0(D5_31), .d1(D13_31), .d2(D21_31), .d3(D29_31),
		.sl0(n27), .sl1(n41) );
	mux4_3 U336 ( .x(n303), .d0(D3_0), .d1(D11_0), .d2(D19_0), .d3(D27_0),
		.sl0(n12), .sl1(n42) );
	mux4_3 U337 ( .x(n304), .d0(D3_1), .d1(D11_1), .d2(D19_1), .d3(D27_1),
		.sl0(n27), .sl1(n42) );
	mux4_3 U338 ( .x(n305), .d0(D3_2), .d1(D11_2), .d2(D19_2), .d3(D27_2),
		.sl0(n27), .sl1(n42) );
	mux4_3 U339 ( .x(n306), .d0(D3_3), .d1(D11_3), .d2(D19_3), .d3(D27_3),
		.sl0(n27), .sl1(n42) );
	mux4_2 U34 ( .x(n237), .d0(n269), .d1(n333), .d2(n301), .d3(n365), .sl0(n10),
		.sl1(n1) );
	mux4_3 U340 ( .x(n307), .d0(D3_4), .d1(D11_4), .d2(D19_4), .d3(D27_4),
		.sl0(n12), .sl1(n42) );
	mux4_3 U341 ( .x(n308), .d0(D3_5), .d1(D11_5), .d2(D19_5), .d3(D27_5),
		.sl0(n21), .sl1(n42) );
	mux4_3 U342 ( .x(n309), .d0(D3_6), .d1(D11_6), .d2(D19_6), .d3(D27_6),
		.sl0(n27), .sl1(n42) );
	mux4_3 U343 ( .x(n310), .d0(D3_7), .d1(D11_7), .d2(D19_7), .d3(D27_7),
		.sl0(n12), .sl1(n42) );
	mux4_3 U344 ( .x(n312), .d0(D3_9), .d1(D11_9), .d2(D19_9), .d3(D27_9),
		.sl0(n21), .sl1(n42) );
	mux4_3 U345 ( .x(n313), .d0(D3_10), .d1(D11_10), .d2(D19_10), .d3(D27_10),
		.sl0(n12), .sl1(n42) );
	mux4_3 U346 ( .x(n314), .d0(D3_11), .d1(D11_11), .d2(D19_11), .d3(D27_11),
		.sl0(n12), .sl1(n42) );
	mux4_3 U347 ( .x(n315), .d0(D3_12), .d1(D11_12), .d2(D19_12), .d3(D27_12),
		.sl0(n12), .sl1(n42) );
	mux4_3 U348 ( .x(n316), .d0(D3_13), .d1(D11_13), .d2(D19_13), .d3(D27_13),
		.sl0(n16), .sl1(n42) );
	mux4_3 U349 ( .x(n317), .d0(D3_14), .d1(D11_14), .d2(D19_14), .d3(D27_14),
		.sl0(n12), .sl1(n42) );
	mux4_2 U35 ( .x(n77), .d0(n109), .d1(n173), .d2(n141), .d3(n205), .sl0(n10),
		.sl1(n1) );
	mux4_3 U350 ( .x(n318), .d0(D3_15), .d1(D11_15), .d2(D19_15), .d3(D27_15),
		.sl0(n13), .sl1(n42) );
	mux4_3 U351 ( .x(n319), .d0(D3_16), .d1(D11_16), .d2(D19_16), .d3(D27_16),
		.sl0(n16), .sl1(n43) );
	mux4_3 U352 ( .x(n320), .d0(D3_17), .d1(D11_17), .d2(D19_17), .d3(D27_17),
		.sl0(n21), .sl1(n43) );
	mux4_3 U353 ( .x(n321), .d0(D3_18), .d1(D11_18), .d2(D19_18), .d3(D27_18),
		.sl0(n21), .sl1(n43) );
	mux4_3 U354 ( .x(n322), .d0(D3_19), .d1(D11_19), .d2(D19_19), .d3(D27_19),
		.sl0(n22), .sl1(n43) );
	mux4_3 U355 ( .x(n323), .d0(D3_20), .d1(D11_20), .d2(D19_20), .d3(D27_20),
		.sl0(n22), .sl1(n43) );
	mux4_3 U356 ( .x(n324), .d0(D3_21), .d1(D11_21), .d2(D19_21), .d3(D27_21),
		.sl0(n22), .sl1(n43) );
	mux4_3 U357 ( .x(n325), .d0(D3_22), .d1(D11_22), .d2(D19_22), .d3(D27_22),
		.sl0(n16), .sl1(n43) );
	mux4_3 U358 ( .x(n326), .d0(D3_23), .d1(D11_23), .d2(D19_23), .d3(D27_23),
		.sl0(n28), .sl1(n43) );
	mux4_3 U359 ( .x(n327), .d0(D3_24), .d1(D11_24), .d2(D19_24), .d3(D27_24),
		.sl0(n22), .sl1(n43) );
	buf_10 U36 ( .x(n1), .a(S2) );
	mux4_3 U360 ( .x(n328), .d0(D3_25), .d1(D11_25), .d2(D19_25), .d3(D27_25),
		.sl0(n26), .sl1(n43) );
	mux4_3 U361 ( .x(n329), .d0(D3_26), .d1(D11_26), .d2(D19_26), .d3(D27_26),
		.sl0(n11), .sl1(n43) );
	mux4_3 U362 ( .x(n330), .d0(D3_27), .d1(D11_27), .d2(D19_27), .d3(D27_27),
		.sl0(n18), .sl1(n43) );
	mux4_3 U363 ( .x(n331), .d0(D3_28), .d1(D11_28), .d2(D19_28), .d3(D27_28),
		.sl0(n11), .sl1(n43) );
	mux4_3 U364 ( .x(n332), .d0(D3_29), .d1(D11_29), .d2(D19_29), .d3(D27_29),
		.sl0(n20), .sl1(n43) );
	mux4_3 U365 ( .x(n333), .d0(D3_30), .d1(D11_30), .d2(D19_30), .d3(D27_30),
		.sl0(n18), .sl1(n43) );
	mux4_3 U366 ( .x(n334), .d0(D3_31), .d1(D11_31), .d2(D19_31), .d3(D27_31),
		.sl0(n20), .sl1(n43) );
	mux4_3 U367 ( .x(n335), .d0(D7_0), .d1(D15_0), .d2(D23_0), .d3(D31_0),
		.sl0(n22), .sl1(n44) );
	mux4_3 U368 ( .x(n336), .d0(D7_1), .d1(D15_1), .d2(D23_1), .d3(D31_1),
		.sl0(n29), .sl1(n44) );
	mux4_3 U369 ( .x(n337), .d0(D7_2), .d1(D15_2), .d2(D23_2), .d3(D31_2),
		.sl0(n22), .sl1(n44) );
	buf_7 U37 ( .x(n2), .a(S2) );
	mux4_3 U370 ( .x(n338), .d0(D7_3), .d1(D15_3), .d2(D23_3), .d3(D31_3),
		.sl0(n28), .sl1(n44) );
	mux4_3 U371 ( .x(n339), .d0(D7_4), .d1(D15_4), .d2(D23_4), .d3(D31_4),
		.sl0(n22), .sl1(n44) );
	mux4_3 U372 ( .x(n340), .d0(D7_5), .d1(D15_5), .d2(D23_5), .d3(D31_5),
		.sl0(n16), .sl1(n44) );
	mux4_3 U373 ( .x(n341), .d0(D7_6), .d1(D15_6), .d2(D23_6), .d3(D31_6),
		.sl0(n11), .sl1(n44) );
	mux4_3 U374 ( .x(n342), .d0(D7_7), .d1(D15_7), .d2(D23_7), .d3(D31_7),
		.sl0(n22), .sl1(n44) );
	mux4_3 U375 ( .x(n343), .d0(D7_8), .d1(D15_8), .d2(D23_8), .d3(D31_8),
		.sl0(n29), .sl1(n44) );
	mux4_3 U376 ( .x(n344), .d0(D7_9), .d1(D15_9), .d2(D23_9), .d3(D31_9),
		.sl0(n22), .sl1(n44) );
	mux4_3 U377 ( .x(n345), .d0(D7_10), .d1(D15_10), .d2(D23_10), .d3(D31_10),
		.sl0(n22), .sl1(n44) );
	mux4_3 U378 ( .x(n346), .d0(D7_11), .d1(D15_11), .d2(D23_11), .d3(D31_11),
		.sl0(n16), .sl1(n44) );
	mux4_3 U379 ( .x(n347), .d0(D7_12), .d1(D15_12), .d2(D23_12), .d3(D31_12),
		.sl0(n26), .sl1(n44) );
	mux4_3 U380 ( .x(n348), .d0(D7_13), .d1(D15_13), .d2(D23_13), .d3(D31_13),
		.sl0(n18), .sl1(n44) );
	mux4_3 U381 ( .x(n349), .d0(D7_14), .d1(D15_14), .d2(D23_14), .d3(D31_14),
		.sl0(n17), .sl1(n44) );
	mux4_3 U382 ( .x(n350), .d0(D7_15), .d1(D15_15), .d2(D23_15), .d3(D31_15),
		.sl0(n22), .sl1(n44) );
	mux4_3 U383 ( .x(n351), .d0(D7_16), .d1(D15_16), .d2(D23_16), .d3(D31_16),
		.sl0(n17), .sl1(n45) );
	mux4_3 U384 ( .x(n352), .d0(D7_17), .d1(D15_17), .d2(D23_17), .d3(D31_17),
		.sl0(n22), .sl1(n45) );
	mux4_3 U385 ( .x(n353), .d0(D7_18), .d1(D15_18), .d2(D23_18), .d3(D31_18),
		.sl0(n20), .sl1(n45) );
	mux4_3 U386 ( .x(n354), .d0(D7_19), .d1(D15_19), .d2(D23_19), .d3(D31_19),
		.sl0(n22), .sl1(n45) );
	mux4_3 U387 ( .x(n355), .d0(D7_20), .d1(D15_20), .d2(D23_20), .d3(D31_20),
		.sl0(n13), .sl1(n45) );
	mux4_3 U388 ( .x(n356), .d0(D7_21), .d1(D15_21), .d2(D23_21), .d3(D31_21),
		.sl0(n13), .sl1(n45) );
	mux4_3 U389 ( .x(n357), .d0(D7_22), .d1(D15_22), .d2(D23_22), .d3(D31_22),
		.sl0(n19), .sl1(n45) );
	buf_14 U39 ( .x(n16), .a(n46) );
	mux4_3 U390 ( .x(n358), .d0(D7_23), .d1(D15_23), .d2(D23_23), .d3(D31_23),
		.sl0(n13), .sl1(n45) );
	mux4_3 U391 ( .x(n359), .d0(D7_24), .d1(D15_24), .d2(D23_24), .d3(D31_24),
		.sl0(n23), .sl1(n45) );
	mux4_3 U392 ( .x(n360), .d0(D7_25), .d1(D15_25), .d2(D23_25), .d3(D31_25),
		.sl0(n23), .sl1(n45) );
	mux4_3 U393 ( .x(n361), .d0(D7_26), .d1(D15_26), .d2(D23_26), .d3(D31_26),
		.sl0(n17), .sl1(n45) );
	mux4_3 U394 ( .x(n362), .d0(D7_27), .d1(D15_27), .d2(D23_27), .d3(D31_27),
		.sl0(n18), .sl1(n45) );
	mux4_3 U395 ( .x(n363), .d0(D7_28), .d1(D15_28), .d2(D23_28), .d3(D31_28),
		.sl0(n16), .sl1(n45) );
	mux4_3 U396 ( .x(n364), .d0(D7_29), .d1(D15_29), .d2(D23_29), .d3(D31_29),
		.sl0(n16), .sl1(n45) );
	mux4_3 U397 ( .x(n365), .d0(D7_30), .d1(D15_30), .d2(D23_30), .d3(D31_30),
		.sl0(n26), .sl1(n45) );
	mux4_3 U398 ( .x(n366), .d0(D7_31), .d1(D15_31), .d2(D23_31), .d3(D31_31),
		.sl0(n11), .sl1(n45) );
	mux2_3 U399 ( .x(Z_0), .d0(n47), .sl(S0), .d1(n207) );
	mux4_2 U4 ( .x(n279), .d0(D5_8), .d1(D13_8), .d2(D21_8), .d3(D29_8), .sl0(n19),
		.sl1(n40) );
	buf_12 U40 ( .x(n28), .a(n46) );
	buf_14 U400 ( .x(n19), .a(n46) );
	inv_16 U401 ( .x(n7), .a(S3) );
	mux2_4 U402 ( .x(Z_25), .d0(n72), .sl(S0), .d1(n232) );
	buf_14 U41 ( .x(n42), .a(S4) );
	buf_10 U42 ( .x(n36), .a(S4) );
	buf_14 U43 ( .x(n37), .a(S4) );
	buf_10 U44 ( .x(n34), .a(S4) );
	buf_10 U45 ( .x(n30), .a(S4) );
	buf_10 U46 ( .x(n40), .a(S4) );
	buf_14 U47 ( .x(n31), .a(S4) );
	buf_12 U48 ( .x(n32), .a(S4) );
	buf_10 U49 ( .x(n33), .a(S4) );
	mux4_2 U5 ( .x(n311), .d0(D3_8), .d1(D11_8), .d2(D19_8), .d3(D27_8), .sl0(n21),
		.sl1(n42) );
	mux4_3 U50 ( .x(n208), .d0(n240), .d1(n304), .d2(n272), .d3(n336), .sl0(S1),
		.sl1(n1) );
	buf_16 U51 ( .x(n4), .a(S1) );
	buf_16 U52 ( .x(n3), .a(S1) );
	buf_10 U53 ( .x(n10), .a(S1) );
	mux2i_3 U54 ( .x(n5), .d0(n208), .sl(n6), .d1(n48) );
	inv_2 U55 ( .x(n6), .a(S0) );
	inv_16 U56 ( .x(n8), .a(n7) );
	buf_10 U57 ( .x(n9), .a(S1) );
	buf_16 U58 ( .x(n11), .a(n46) );
	buf_16 U59 ( .x(n12), .a(n8) );
	mux4_2 U6 ( .x(n183), .d0(D6_8), .d1(D14_8), .d2(D22_8), .d3(D30_8), .sl0(n14),
		.sl1(n36) );
	buf_16 U60 ( .x(n13), .a(n46) );
	buf_16 U61 ( .x(n14), .a(n8) );
	buf_16 U62 ( .x(n15), .a(n8) );
	buf_16 U63 ( .x(n17), .a(n46) );
	buf_16 U64 ( .x(n18), .a(n46) );
	buf_16 U66 ( .x(n20), .a(n46) );
	buf_16 U67 ( .x(n21), .a(n8) );
	buf_16 U68 ( .x(n22), .a(n8) );
	buf_16 U69 ( .x(n23), .a(n8) );
	mux4_2 U7 ( .x(n119), .d0(D4_8), .d1(D12_8), .d2(D20_8), .d3(D28_8), .sl0(n24),
		.sl1(n32) );
	buf_16 U70 ( .x(n24), .a(n8) );
	buf_16 U71 ( .x(n25), .a(n8) );
	buf_16 U72 ( .x(n26), .a(n46) );
	buf_16 U73 ( .x(n27), .a(n8) );
	buf_16 U74 ( .x(n29), .a(n46) );
	buf_16 U75 ( .x(n38), .a(S4) );
	buf_16 U76 ( .x(n39), .a(S4) );
	buf_16 U77 ( .x(n43), .a(S4) );
	buf_16 U78 ( .x(n44), .a(S4) );
	buf_16 U79 ( .x(n45), .a(S4) );
	mux4_2 U8 ( .x(n87), .d0(D0_8), .d1(D8_8), .d2(D16_8), .d3(D24_8), .sl0(n23),
		.sl1(n30) );
	inv_16 U80 ( .x(n46), .a(n7) );
	mux2_4 U82 ( .x(Z_2), .d0(n49), .sl(S0), .d1(n209) );
	mux2_4 U83 ( .x(Z_3), .d0(n50), .sl(S0), .d1(n210) );
	mux2_4 U84 ( .x(Z_4), .d0(n51), .sl(S0), .d1(n211) );
	mux2_4 U85 ( .x(Z_5), .d0(n52), .sl(S0), .d1(n212) );
	mux2_4 U86 ( .x(Z_6), .d0(n53), .sl(S0), .d1(n213) );
	mux2_4 U87 ( .x(Z_7), .d0(n54), .sl(S0), .d1(n214) );
	mux2_4 U88 ( .x(Z_8), .d0(n55), .sl(S0), .d1(n215) );
	mux2_4 U89 ( .x(Z_9), .d0(n56), .sl(S0), .d1(n216) );
	mux4_2 U9 ( .x(n282), .d0(D5_11), .d1(D13_11), .d2(D21_11), .d3(D29_11),
		.sl0(n12), .sl1(n40) );
	mux2_4 U90 ( .x(Z_10), .d0(n57), .sl(S0), .d1(n217) );
	mux2_4 U91 ( .x(Z_11), .d0(n58), .sl(S0), .d1(n218) );
	mux2_4 U92 ( .x(Z_12), .d0(n59), .sl(S0), .d1(n219) );
	mux2_4 U93 ( .x(Z_13), .d0(n60), .sl(S0), .d1(n220) );
	mux2_4 U94 ( .x(Z_14), .d0(n61), .sl(S0), .d1(n221) );
	mux2_4 U95 ( .x(Z_15), .d0(n62), .sl(S0), .d1(n222) );
	mux2_4 U96 ( .x(Z_16), .d0(n63), .sl(S0), .d1(n223) );
	mux2_4 U97 ( .x(Z_17), .d0(n64), .sl(S0), .d1(n224) );
	mux2_4 U98 ( .x(Z_18), .d0(n65), .sl(S0), .d1(n225) );
	mux2_4 U99 ( .x(Z_19), .d0(n66), .sl(S0), .d1(n226) );

endmodule


module DLX_sync_MUX_OP_32_5_32_test_1 (  D0_31, D0_30, D0_29, D0_28, D0_27,
	D0_26, D0_25, D0_24, D0_23, D0_22, D0_21, D0_20, D0_19, D0_18, D0_17,
	D0_16, D0_15, D0_14, D0_13, D0_12, D0_11, D0_10, D0_9, D0_8, D0_7, D0_6,
	D0_5, D0_4, D0_3, D0_2, D0_1, D0_0, D1_31, D1_30, D1_29, D1_28, D1_27,
	D1_26, D1_25, D1_24, D1_23, D1_22, D1_21, D1_20, D1_19, D1_18, D1_17,
	D1_16, D1_15, D1_14, D1_13, D1_12, D1_11, D1_10, D1_9, D1_8, D1_7, D1_6,
	D1_5, D1_4, D1_3, D1_2, D1_1, D1_0, D2_31, D2_30, D2_29, D2_28, D2_27,
	D2_26, D2_25, D2_24, D2_23, D2_22, D2_21, D2_20, D2_19, D2_18, D2_17,
	D2_16, D2_15, D2_14, D2_13, D2_12, D2_11, D2_10, D2_9, D2_8, D2_7, D2_6,
	D2_5, D2_4, D2_3, D2_2, D2_1, D2_0, D3_31, D3_30, D3_29, D3_28, D3_27,
	D3_26, D3_25, D3_24, D3_23, D3_22, D3_21, D3_20, D3_19, D3_18, D3_17,
	D3_16, D3_15, D3_14, D3_13, D3_12, D3_11, D3_10, D3_9, D3_8, D3_7, D3_6,
	D3_5, D3_4, D3_3, D3_2, D3_1, D3_0, D4_31, D4_30, D4_29, D4_28, D4_27,
	D4_26, D4_25, D4_24, D4_23, D4_22, D4_21, D4_20, D4_19, D4_18, D4_17,
	D4_16, D4_15, D4_14, D4_13, D4_12, D4_11, D4_10, D4_9, D4_8, D4_7, D4_6,
	D4_5, D4_4, D4_3, D4_2, D4_1, D4_0, D5_31, D5_30, D5_29, D5_28, D5_27,
	D5_26, D5_25, D5_24, D5_23, D5_22, D5_21, D5_20, D5_19, D5_18, D5_17,
	D5_16, D5_15, D5_14, D5_13, D5_12, D5_11, D5_10, D5_9, D5_8, D5_7, D5_6,
	D5_5, D5_4, D5_3, D5_2, D5_1, D5_0, D6_31, D6_30, D6_29, D6_28, D6_27,
	D6_26, D6_25, D6_24, D6_23, D6_22, D6_21, D6_20, D6_19, D6_18, D6_17,
	D6_16, D6_15, D6_14, D6_13, D6_12, D6_11, D6_10, D6_9, D6_8, D6_7, D6_6,
	D6_5, D6_4, D6_3, D6_2, D6_1, D6_0, D7_31, D7_30, D7_29, D7_28, D7_27,
	D7_26, D7_25, D7_24, D7_23, D7_22, D7_21, D7_20, D7_19, D7_18, D7_17,
	D7_16, D7_15, D7_14, D7_13, D7_12, D7_11, D7_10, D7_9, D7_8, D7_7, D7_6,
	D7_5, D7_4, D7_3, D7_2, D7_1, D7_0, D8_31, D8_30, D8_29, D8_28, D8_27,
	D8_26, D8_25, D8_24, D8_23, D8_22, D8_21, D8_20, D8_19, D8_18, D8_17,
	D8_16, D8_15, D8_14, D8_13, D8_12, D8_11, D8_10, D8_9, D8_8, D8_7, D8_6,
	D8_5, D8_4, D8_3, D8_2, D8_1, D8_0, D9_31, D9_30, D9_29, D9_28, D9_27,
	D9_26, D9_25, D9_24, D9_23, D9_22, D9_21, D9_20, D9_19, D9_18, D9_17,
	D9_16, D9_15, D9_14, D9_13, D9_12, D9_11, D9_10, D9_9, D9_8, D9_7, D9_6,
	D9_5, D9_4, D9_3, D9_2, D9_1, D9_0, D10_31, D10_30, D10_29, D10_28, D10_27,
	D10_26, D10_25, D10_24, D10_23, D10_22, D10_21, D10_20, D10_19, D10_18,
	D10_17, D10_16, D10_15, D10_14, D10_13, D10_12, D10_11, D10_10, D10_9,
	D10_8, D10_7, D10_6, D10_5, D10_4, D10_3, D10_2, D10_1, D10_0, D11_31,
	D11_30, D11_29, D11_28, D11_27, D11_26, D11_25, D11_24, D11_23, D11_22,
	D11_21, D11_20, D11_19, D11_18, D11_17, D11_16, D11_15, D11_14, D11_13,
	D11_12, D11_11, D11_10, D11_9, D11_8, D11_7, D11_6, D11_5, D11_4, D11_3,
	D11_2, D11_1, D11_0, D12_31, D12_30, D12_29, D12_28, D12_27, D12_26, D12_25,
	D12_24, D12_23, D12_22, D12_21, D12_20, D12_19, D12_18, D12_17, D12_16,
	D12_15, D12_14, D12_13, D12_12, D12_11, D12_10, D12_9, D12_8, D12_7, D12_6,
	D12_5, D12_4, D12_3, D12_2, D12_1, D12_0, D13_31, D13_30, D13_29, D13_28,
	D13_27, D13_26, D13_25, D13_24, D13_23, D13_22, D13_21, D13_20, D13_19,
	D13_18, D13_17, D13_16, D13_15, D13_14, D13_13, D13_12, D13_11, D13_10,
	D13_9, D13_8, D13_7, D13_6, D13_5, D13_4, D13_3, D13_2, D13_1, D13_0,
	D14_31, D14_30, D14_29, D14_28, D14_27, D14_26, D14_25, D14_24, D14_23,
	D14_22, D14_21, D14_20, D14_19, D14_18, D14_17, D14_16, D14_15, D14_14,
	D14_13, D14_12, D14_11, D14_10, D14_9, D14_8, D14_7, D14_6, D14_5, D14_4,
	D14_3, D14_2, D14_1, D14_0, D15_31, D15_30, D15_29, D15_28, D15_27, D15_26,
	D15_25, D15_24, D15_23, D15_22, D15_21, D15_20, D15_19, D15_18, D15_17,
	D15_16, D15_15, D15_14, D15_13, D15_12, D15_11, D15_10, D15_9, D15_8,
	D15_7, D15_6, D15_5, D15_4, D15_3, D15_2, D15_1, D15_0, D16_31, D16_30,
	D16_29, D16_28, D16_27, D16_26, D16_25, D16_24, D16_23, D16_22, D16_21,
	D16_20, D16_19, D16_18, D16_17, D16_16, D16_15, D16_14, D16_13, D16_12,
	D16_11, D16_10, D16_9, D16_8, D16_7, D16_6, D16_5, D16_4, D16_3, D16_2,
	D16_1, D16_0, D17_31, D17_30, D17_29, D17_28, D17_27, D17_26, D17_25,
	D17_24, D17_23, D17_22, D17_21, D17_20, D17_19, D17_18, D17_17, D17_16,
	D17_15, D17_14, D17_13, D17_12, D17_11, D17_10, D17_9, D17_8, D17_7, D17_6,
	D17_5, D17_4, D17_3, D17_2, D17_1, D17_0, D18_31, D18_30, D18_29, D18_28,
	D18_27, D18_26, D18_25, D18_24, D18_23, D18_22, D18_21, D18_20, D18_19,
	D18_18, D18_17, D18_16, D18_15, D18_14, D18_13, D18_12, D18_11, D18_10,
	D18_9, D18_8, D18_7, D18_6, D18_5, D18_4, D18_3, D18_2, D18_1, D18_0,
	D19_31, D19_30, D19_29, D19_28, D19_27, D19_26, D19_25, D19_24, D19_23,
	D19_22, D19_21, D19_20, D19_19, D19_18, D19_17, D19_16, D19_15, D19_14,
	D19_13, D19_12, D19_11, D19_10, D19_9, D19_8, D19_7, D19_6, D19_5, D19_4,
	D19_3, D19_2, D19_1, D19_0, D20_31, D20_30, D20_29, D20_28, D20_27, D20_26,
	D20_25, D20_24, D20_23, D20_22, D20_21, D20_20, D20_19, D20_18, D20_17,
	D20_16, D20_15, D20_14, D20_13, D20_12, D20_11, D20_10, D20_9, D20_8,
	D20_7, D20_6, D20_5, D20_4, D20_3, D20_2, D20_1, D20_0, D21_31, D21_30,
	D21_29, D21_28, D21_27, D21_26, D21_25, D21_24, D21_23, D21_22, D21_21,
	D21_20, D21_19, D21_18, D21_17, D21_16, D21_15, D21_14, D21_13, D21_12,
	D21_11, D21_10, D21_9, D21_8, D21_7, D21_6, D21_5, D21_4, D21_3, D21_2,
	D21_1, D21_0, D22_31, D22_30, D22_29, D22_28, D22_27, D22_26, D22_25,
	D22_24, D22_23, D22_22, D22_21, D22_20, D22_19, D22_18, D22_17, D22_16,
	D22_15, D22_14, D22_13, D22_12, D22_11, D22_10, D22_9, D22_8, D22_7, D22_6,
	D22_5, D22_4, D22_3, D22_2, D22_1, D22_0, D23_31, D23_30, D23_29, D23_28,
	D23_27, D23_26, D23_25, D23_24, D23_23, D23_22, D23_21, D23_20, D23_19,
	D23_18, D23_17, D23_16, D23_15, D23_14, D23_13, D23_12, D23_11, D23_10,
	D23_9, D23_8, D23_7, D23_6, D23_5, D23_4, D23_3, D23_2, D23_1, D23_0,
	D24_31, D24_30, D24_29, D24_28, D24_27, D24_26, D24_25, D24_24, D24_23,
	D24_22, D24_21, D24_20, D24_19, D24_18, D24_17, D24_16, D24_15, D24_14,
	D24_13, D24_12, D24_11, D24_10, D24_9, D24_8, D24_7, D24_6, D24_5, D24_4,
	D24_3, D24_2, D24_1, D24_0, D25_31, D25_30, D25_29, D25_28, D25_27, D25_26,
	D25_25, D25_24, D25_23, D25_22, D25_21, D25_20, D25_19, D25_18, D25_17,
	D25_16, D25_15, D25_14, D25_13, D25_12, D25_11, D25_10, D25_9, D25_8,
	D25_7, D25_6, D25_5, D25_4, D25_3, D25_2, D25_1, D25_0, D26_31, D26_30,
	D26_29, D26_28, D26_27, D26_26, D26_25, D26_24, D26_23, D26_22, D26_21,
	D26_20, D26_19, D26_18, D26_17, D26_16, D26_15, D26_14, D26_13, D26_12,
	D26_11, D26_10, D26_9, D26_8, D26_7, D26_6, D26_5, D26_4, D26_3, D26_2,
	D26_1, D26_0, D27_31, D27_30, D27_29, D27_28, D27_27, D27_26, D27_25,
	D27_24, D27_23, D27_22, D27_21, D27_20, D27_19, D27_18, D27_17, D27_16,
	D27_15, D27_14, D27_13, D27_12, D27_11, D27_10, D27_9, D27_8, D27_7, D27_6,
	D27_5, D27_4, D27_3, D27_2, D27_1, D27_0, D28_31, D28_30, D28_29, D28_28,
	D28_27, D28_26, D28_25, D28_24, D28_23, D28_22, D28_21, D28_20, D28_19,
	D28_18, D28_17, D28_16, D28_15, D28_14, D28_13, D28_12, D28_11, D28_10,
	D28_9, D28_8, D28_7, D28_6, D28_5, D28_4, D28_3, D28_2, D28_1, D28_0,
	D29_31, D29_30, D29_29, D29_28, D29_27, D29_26, D29_25, D29_24, D29_23,
	D29_22, D29_21, D29_20, D29_19, D29_18, D29_17, D29_16, D29_15, D29_14,
	D29_13, D29_12, D29_11, D29_10, D29_9, D29_8, D29_7, D29_6, D29_5, D29_4,
	D29_3, D29_2, D29_1, D29_0, D30_31, D30_30, D30_29, D30_28, D30_27, D30_26,
	D30_25, D30_24, D30_23, D30_22, D30_21, D30_20, D30_19, D30_18, D30_17,
	D30_16, D30_15, D30_14, D30_13, D30_12, D30_11, D30_10, D30_9, D30_8,
	D30_7, D30_6, D30_5, D30_4, D30_3, D30_2, D30_1, D30_0, D31_31, D31_30,
	D31_29, D31_28, D31_27, D31_26, D31_25, D31_24, D31_23, D31_22, D31_21,
	D31_20, D31_19, D31_18, D31_17, D31_16, D31_15, D31_14, D31_13, D31_12,
	D31_11, D31_10, D31_9, D31_8, D31_7, D31_6, D31_5, D31_4, D31_3, D31_2,
	D31_1, D31_0, S0, S1, S2, S3, S4, Z_31, Z_30, Z_29, Z_28, Z_27, Z_26,
	Z_25, Z_24, Z_23, Z_22, Z_21, Z_20, Z_19, Z_18, Z_17, Z_16, Z_15, Z_14,
	Z_13, Z_12, Z_11, Z_10, Z_9, Z_8, Z_7, Z_6, Z_5, Z_4, Z_3, Z_2, Z_1, Z_0 );

input  D0_31, D0_30, D0_29, D0_28, D0_27, D0_26, D0_25, D0_24, D0_23, D0_22,
	D0_21, D0_20, D0_19, D0_18, D0_17, D0_16, D0_15, D0_14, D0_13, D0_12,
	D0_11, D0_10, D0_9, D0_8, D0_7, D0_6, D0_5, D0_4, D0_3, D0_2, D0_1, D0_0,
	D1_31, D1_30, D1_29, D1_28, D1_27, D1_26, D1_25, D1_24, D1_23, D1_22,
	D1_21, D1_20, D1_19, D1_18, D1_17, D1_16, D1_15, D1_14, D1_13, D1_12,
	D1_11, D1_10, D1_9, D1_8, D1_7, D1_6, D1_5, D1_4, D1_3, D1_2, D1_1, D1_0,
	D2_31, D2_30, D2_29, D2_28, D2_27, D2_26, D2_25, D2_24, D2_23, D2_22,
	D2_21, D2_20, D2_19, D2_18, D2_17, D2_16, D2_15, D2_14, D2_13, D2_12,
	D2_11, D2_10, D2_9, D2_8, D2_7, D2_6, D2_5, D2_4, D2_3, D2_2, D2_1, D2_0,
	D3_31, D3_30, D3_29, D3_28, D3_27, D3_26, D3_25, D3_24, D3_23, D3_22,
	D3_21, D3_20, D3_19, D3_18, D3_17, D3_16, D3_15, D3_14, D3_13, D3_12,
	D3_11, D3_10, D3_9, D3_8, D3_7, D3_6, D3_5, D3_4, D3_3, D3_2, D3_1, D3_0,
	D4_31, D4_30, D4_29, D4_28, D4_27, D4_26, D4_25, D4_24, D4_23, D4_22,
	D4_21, D4_20, D4_19, D4_18, D4_17, D4_16, D4_15, D4_14, D4_13, D4_12,
	D4_11, D4_10, D4_9, D4_8, D4_7, D4_6, D4_5, D4_4, D4_3, D4_2, D4_1, D4_0,
	D5_31, D5_30, D5_29, D5_28, D5_27, D5_26, D5_25, D5_24, D5_23, D5_22,
	D5_21, D5_20, D5_19, D5_18, D5_17, D5_16, D5_15, D5_14, D5_13, D5_12,
	D5_11, D5_10, D5_9, D5_8, D5_7, D5_6, D5_5, D5_4, D5_3, D5_2, D5_1, D5_0,
	D6_31, D6_30, D6_29, D6_28, D6_27, D6_26, D6_25, D6_24, D6_23, D6_22,
	D6_21, D6_20, D6_19, D6_18, D6_17, D6_16, D6_15, D6_14, D6_13, D6_12,
	D6_11, D6_10, D6_9, D6_8, D6_7, D6_6, D6_5, D6_4, D6_3, D6_2, D6_1, D6_0,
	D7_31, D7_30, D7_29, D7_28, D7_27, D7_26, D7_25, D7_24, D7_23, D7_22,
	D7_21, D7_20, D7_19, D7_18, D7_17, D7_16, D7_15, D7_14, D7_13, D7_12,
	D7_11, D7_10, D7_9, D7_8, D7_7, D7_6, D7_5, D7_4, D7_3, D7_2, D7_1, D7_0,
	D8_31, D8_30, D8_29, D8_28, D8_27, D8_26, D8_25, D8_24, D8_23, D8_22,
	D8_21, D8_20, D8_19, D8_18, D8_17, D8_16, D8_15, D8_14, D8_13, D8_12,
	D8_11, D8_10, D8_9, D8_8, D8_7, D8_6, D8_5, D8_4, D8_3, D8_2, D8_1, D8_0,
	D9_31, D9_30, D9_29, D9_28, D9_27, D9_26, D9_25, D9_24, D9_23, D9_22,
	D9_21, D9_20, D9_19, D9_18, D9_17, D9_16, D9_15, D9_14, D9_13, D9_12,
	D9_11, D9_10, D9_9, D9_8, D9_7, D9_6, D9_5, D9_4, D9_3, D9_2, D9_1, D9_0,
	D10_31, D10_30, D10_29, D10_28, D10_27, D10_26, D10_25, D10_24, D10_23,
	D10_22, D10_21, D10_20, D10_19, D10_18, D10_17, D10_16, D10_15, D10_14,
	D10_13, D10_12, D10_11, D10_10, D10_9, D10_8, D10_7, D10_6, D10_5, D10_4,
	D10_3, D10_2, D10_1, D10_0, D11_31, D11_30, D11_29, D11_28, D11_27, D11_26,
	D11_25, D11_24, D11_23, D11_22, D11_21, D11_20, D11_19, D11_18, D11_17,
	D11_16, D11_15, D11_14, D11_13, D11_12, D11_11, D11_10, D11_9, D11_8,
	D11_7, D11_6, D11_5, D11_4, D11_3, D11_2, D11_1, D11_0, D12_31, D12_30,
	D12_29, D12_28, D12_27, D12_26, D12_25, D12_24, D12_23, D12_22, D12_21,
	D12_20, D12_19, D12_18, D12_17, D12_16, D12_15, D12_14, D12_13, D12_12,
	D12_11, D12_10, D12_9, D12_8, D12_7, D12_6, D12_5, D12_4, D12_3, D12_2,
	D12_1, D12_0, D13_31, D13_30, D13_29, D13_28, D13_27, D13_26, D13_25,
	D13_24, D13_23, D13_22, D13_21, D13_20, D13_19, D13_18, D13_17, D13_16,
	D13_15, D13_14, D13_13, D13_12, D13_11, D13_10, D13_9, D13_8, D13_7, D13_6,
	D13_5, D13_4, D13_3, D13_2, D13_1, D13_0, D14_31, D14_30, D14_29, D14_28,
	D14_27, D14_26, D14_25, D14_24, D14_23, D14_22, D14_21, D14_20, D14_19,
	D14_18, D14_17, D14_16, D14_15, D14_14, D14_13, D14_12, D14_11, D14_10,
	D14_9, D14_8, D14_7, D14_6, D14_5, D14_4, D14_3, D14_2, D14_1, D14_0,
	D15_31, D15_30, D15_29, D15_28, D15_27, D15_26, D15_25, D15_24, D15_23,
	D15_22, D15_21, D15_20, D15_19, D15_18, D15_17, D15_16, D15_15, D15_14,
	D15_13, D15_12, D15_11, D15_10, D15_9, D15_8, D15_7, D15_6, D15_5, D15_4,
	D15_3, D15_2, D15_1, D15_0, D16_31, D16_30, D16_29, D16_28, D16_27, D16_26,
	D16_25, D16_24, D16_23, D16_22, D16_21, D16_20, D16_19, D16_18, D16_17,
	D16_16, D16_15, D16_14, D16_13, D16_12, D16_11, D16_10, D16_9, D16_8,
	D16_7, D16_6, D16_5, D16_4, D16_3, D16_2, D16_1, D16_0, D17_31, D17_30,
	D17_29, D17_28, D17_27, D17_26, D17_25, D17_24, D17_23, D17_22, D17_21,
	D17_20, D17_19, D17_18, D17_17, D17_16, D17_15, D17_14, D17_13, D17_12,
	D17_11, D17_10, D17_9, D17_8, D17_7, D17_6, D17_5, D17_4, D17_3, D17_2,
	D17_1, D17_0, D18_31, D18_30, D18_29, D18_28, D18_27, D18_26, D18_25,
	D18_24, D18_23, D18_22, D18_21, D18_20, D18_19, D18_18, D18_17, D18_16,
	D18_15, D18_14, D18_13, D18_12, D18_11, D18_10, D18_9, D18_8, D18_7, D18_6,
	D18_5, D18_4, D18_3, D18_2, D18_1, D18_0, D19_31, D19_30, D19_29, D19_28,
	D19_27, D19_26, D19_25, D19_24, D19_23, D19_22, D19_21, D19_20, D19_19,
	D19_18, D19_17, D19_16, D19_15, D19_14, D19_13, D19_12, D19_11, D19_10,
	D19_9, D19_8, D19_7, D19_6, D19_5, D19_4, D19_3, D19_2, D19_1, D19_0,
	D20_31, D20_30, D20_29, D20_28, D20_27, D20_26, D20_25, D20_24, D20_23,
	D20_22, D20_21, D20_20, D20_19, D20_18, D20_17, D20_16, D20_15, D20_14,
	D20_13, D20_12, D20_11, D20_10, D20_9, D20_8, D20_7, D20_6, D20_5, D20_4,
	D20_3, D20_2, D20_1, D20_0, D21_31, D21_30, D21_29, D21_28, D21_27, D21_26,
	D21_25, D21_24, D21_23, D21_22, D21_21, D21_20, D21_19, D21_18, D21_17,
	D21_16, D21_15, D21_14, D21_13, D21_12, D21_11, D21_10, D21_9, D21_8,
	D21_7, D21_6, D21_5, D21_4, D21_3, D21_2, D21_1, D21_0, D22_31, D22_30,
	D22_29, D22_28, D22_27, D22_26, D22_25, D22_24, D22_23, D22_22, D22_21,
	D22_20, D22_19, D22_18, D22_17, D22_16, D22_15, D22_14, D22_13, D22_12,
	D22_11, D22_10, D22_9, D22_8, D22_7, D22_6, D22_5, D22_4, D22_3, D22_2,
	D22_1, D22_0, D23_31, D23_30, D23_29, D23_28, D23_27, D23_26, D23_25,
	D23_24, D23_23, D23_22, D23_21, D23_20, D23_19, D23_18, D23_17, D23_16,
	D23_15, D23_14, D23_13, D23_12, D23_11, D23_10, D23_9, D23_8, D23_7, D23_6,
	D23_5, D23_4, D23_3, D23_2, D23_1, D23_0, D24_31, D24_30, D24_29, D24_28,
	D24_27, D24_26, D24_25, D24_24, D24_23, D24_22, D24_21, D24_20, D24_19,
	D24_18, D24_17, D24_16, D24_15, D24_14, D24_13, D24_12, D24_11, D24_10,
	D24_9, D24_8, D24_7, D24_6, D24_5, D24_4, D24_3, D24_2, D24_1, D24_0,
	D25_31, D25_30, D25_29, D25_28, D25_27, D25_26, D25_25, D25_24, D25_23,
	D25_22, D25_21, D25_20, D25_19, D25_18, D25_17, D25_16, D25_15, D25_14,
	D25_13, D25_12, D25_11, D25_10, D25_9, D25_8, D25_7, D25_6, D25_5, D25_4,
	D25_3, D25_2, D25_1, D25_0, D26_31, D26_30, D26_29, D26_28, D26_27, D26_26,
	D26_25, D26_24, D26_23, D26_22, D26_21, D26_20, D26_19, D26_18, D26_17,
	D26_16, D26_15, D26_14, D26_13, D26_12, D26_11, D26_10, D26_9, D26_8,
	D26_7, D26_6, D26_5, D26_4, D26_3, D26_2, D26_1, D26_0, D27_31, D27_30,
	D27_29, D27_28, D27_27, D27_26, D27_25, D27_24, D27_23, D27_22, D27_21,
	D27_20, D27_19, D27_18, D27_17, D27_16, D27_15, D27_14, D27_13, D27_12,
	D27_11, D27_10, D27_9, D27_8, D27_7, D27_6, D27_5, D27_4, D27_3, D27_2,
	D27_1, D27_0, D28_31, D28_30, D28_29, D28_28, D28_27, D28_26, D28_25,
	D28_24, D28_23, D28_22, D28_21, D28_20, D28_19, D28_18, D28_17, D28_16,
	D28_15, D28_14, D28_13, D28_12, D28_11, D28_10, D28_9, D28_8, D28_7, D28_6,
	D28_5, D28_4, D28_3, D28_2, D28_1, D28_0, D29_31, D29_30, D29_29, D29_28,
	D29_27, D29_26, D29_25, D29_24, D29_23, D29_22, D29_21, D29_20, D29_19,
	D29_18, D29_17, D29_16, D29_15, D29_14, D29_13, D29_12, D29_11, D29_10,
	D29_9, D29_8, D29_7, D29_6, D29_5, D29_4, D29_3, D29_2, D29_1, D29_0,
	D30_31, D30_30, D30_29, D30_28, D30_27, D30_26, D30_25, D30_24, D30_23,
	D30_22, D30_21, D30_20, D30_19, D30_18, D30_17, D30_16, D30_15, D30_14,
	D30_13, D30_12, D30_11, D30_10, D30_9, D30_8, D30_7, D30_6, D30_5, D30_4,
	D30_3, D30_2, D30_1, D30_0, D31_31, D31_30, D31_29, D31_28, D31_27, D31_26,
	D31_25, D31_24, D31_23, D31_22, D31_21, D31_20, D31_19, D31_18, D31_17,
	D31_16, D31_15, D31_14, D31_13, D31_12, D31_11, D31_10, D31_9, D31_8,
	D31_7, D31_6, D31_5, D31_4, D31_3, D31_2, D31_1, D31_0, S0, S1, S2, S3,
	S4;
output  Z_31, Z_30, Z_29, Z_28, Z_27, Z_26, Z_25, Z_24, Z_23, Z_22, Z_21,
	Z_20, Z_19, Z_18, Z_17, Z_16, Z_15, Z_14, Z_13, Z_12, Z_11, Z_10, Z_9,
	Z_8, Z_7, Z_6, Z_5, Z_4, Z_3, Z_2, Z_1, Z_0;

wire n1, n10, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
	n11, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n12,
	n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n13, n130,
	n131, n132, n133, n134, n135, n136, n137, n138, n139, n14, n140, n141,
	n142, n1425, n143, n144, n145, n146, n147, n148, n149, n15, n150, n151,
	n152, n153, n154, n155, n156, n157, n158, n159, n16, n160, n161, n162,
	n163, n164, n165, n166, n167, n168, n169, n17, n170, n171, n172, n173,
	n174, n175, n176, n177, n178, n179, n18, n180, n181, n182, n183, n184,
	n185, n186, n187, n188, n189, n19, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n2, n20, n200, n201, n202, n203, n204, n205, n206,
	n207, n208, n209, n21, n210, n211, n212, n213, n214, n215, n216, n217,
	n218, n219, n22, n220, n221, n222, n223, n224, n225, n226, n227, n228,
	n229, n23, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
	n24, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n25,
	n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n26, n260,
	n261, n262, n263, n264, n265, n266, n267, n268, n269, n27, n270, n271,
	n272, n273, n274, n275, n276, n277, n278, n279, n28, n280, n281, n282,
	n283, n284, n285, n286, n287, n288, n289, n29, n290, n291, n292, n293,
	n294, n295, n296, n297, n298, n299, n3, n30, n300, n301, n302, n303, n304,
	n305, n306, n307, n308, n309, n31, n310, n311, n312, n313, n314, n315,
	n316, n317, n318, n319, n32, n320, n321, n322, n323, n324, n325, n326,
	n327, n328, n329, n33, n330, n331, n332, n333, n334, n335, n336, n337,
	n338, n339, n34, n340, n341, n342, n343, n344, n345, n346, n347, n348,
	n349, n35, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
	n36, n360, n361, n362, n363, n37, n38, n39, n4, n40, n41, n42, n43, n44,
	n45, n46, n47, n48, n49, n5, n50, n51, n52, n53, n54, n55, n56, n57, n58,
	n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n7, n70, n71, n72,
	n73, n74, n75, n76, n77, n78, n79, n8, n80, n81, n82, n83, n84, n85, n86,
	n87, n88, n89, n9, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	mux4_1 U1 ( .x(n342), .d0(D7_10), .d1(D15_10), .d2(D23_10), .d3(D31_10),
		.sl0(n18), .sl1(n40) );
	mux4_1 U10 ( .x(n299), .d0(D5_31), .d1(D13_31), .d2(D21_31), .d3(D29_31),
		.sl0(n8), .sl1(n37) );
	mux4_1 U100 ( .x(n249), .d0(D1_13), .d1(D9_13), .d2(D17_13), .d3(D25_13),
		.sl0(n22), .sl1(n34) );
	mux4_1 U101 ( .x(n185), .d0(D6_13), .d1(D14_13), .d2(D22_13), .d3(D30_13),
		.sl0(n15), .sl1(n32) );
	mux4_1 U102 ( .x(n121), .d0(D4_13), .d1(D12_13), .d2(D20_13), .d3(D28_13),
		.sl0(n11), .sl1(n28) );
	mux4_1 U103 ( .x(n153), .d0(D2_13), .d1(D10_13), .d2(D18_13), .d3(D26_13),
		.sl0(n20), .sl1(n30) );
	mux4_1 U104 ( .x(n89), .d0(D0_13), .d1(D8_13), .d2(D16_13), .d3(D24_13),
		.sl0(n19), .sl1(n26) );
	mux4_1 U105 ( .x(n350), .d0(D7_18), .d1(D15_18), .d2(D23_18), .d3(D31_18),
		.sl0(n24), .sl1(n41) );
	mux4_1 U106 ( .x(n286), .d0(D5_18), .d1(D13_18), .d2(D21_18), .d3(D29_18),
		.sl0(n23), .sl1(n37) );
	mux4_1 U107 ( .x(n318), .d0(D3_18), .d1(D11_18), .d2(D19_18), .d3(D27_18),
		.sl0(n18), .sl1(n39) );
	mux4_1 U108 ( .x(n254), .d0(D1_18), .d1(D9_18), .d2(D17_18), .d3(D25_18),
		.sl0(n22), .sl1(n35) );
	mux4_1 U109 ( .x(n190), .d0(D6_18), .d1(D14_18), .d2(D22_18), .d3(D30_18),
		.sl0(n21), .sl1(n33) );
	mux4_1 U11 ( .x(n331), .d0(D3_31), .d1(D11_31), .d2(D19_31), .d3(D27_31),
		.sl0(n18), .sl1(n39) );
	mux4_1 U110 ( .x(n126), .d0(D4_18), .d1(D12_18), .d2(D20_18), .d3(D28_18),
		.sl0(n20), .sl1(n29) );
	mux4_1 U111 ( .x(n158), .d0(D2_18), .d1(D10_18), .d2(D18_18), .d3(D26_18),
		.sl0(n11), .sl1(n31) );
	mux4_1 U112 ( .x(n94), .d0(D0_18), .d1(D8_18), .d2(D16_18), .d3(D24_18),
		.sl0(n19), .sl1(n27) );
	mux4_1 U113 ( .x(n344), .d0(D7_12), .d1(D15_12), .d2(D23_12), .d3(D31_12),
		.sl0(n7), .sl1(n40) );
	mux4_1 U114 ( .x(n280), .d0(D5_12), .d1(D13_12), .d2(D21_12), .d3(D29_12),
		.sl0(n8), .sl1(n36) );
	mux4_1 U115 ( .x(n312), .d0(D3_12), .d1(D11_12), .d2(D19_12), .d3(D27_12),
		.sl0(n8), .sl1(n38) );
	mux4_1 U116 ( .x(n248), .d0(D1_12), .d1(D9_12), .d2(D17_12), .d3(D25_12),
		.sl0(n16), .sl1(n34) );
	mux4_1 U117 ( .x(n184), .d0(D6_12), .d1(D14_12), .d2(D22_12), .d3(D30_12),
		.sl0(n15), .sl1(n32) );
	mux4_1 U118 ( .x(n120), .d0(D4_12), .d1(D12_12), .d2(D20_12), .d3(D28_12),
		.sl0(n20), .sl1(n28) );
	mux4_1 U119 ( .x(n152), .d0(D2_12), .d1(D10_12), .d2(D18_12), .d3(D26_12),
		.sl0(n20), .sl1(n30) );
	mux4_1 U12 ( .x(n267), .d0(D1_31), .d1(D9_31), .d2(D17_31), .d3(D25_31),
		.sl0(n9), .sl1(n35) );
	mux4_1 U120 ( .x(n88), .d0(D0_12), .d1(D8_12), .d2(D16_12), .d3(D24_12),
		.sl0(n13), .sl1(n26) );
	mux4_1 U121 ( .x(n349), .d0(D7_17), .d1(D15_17), .d2(D23_17), .d3(D31_17),
		.sl0(n18), .sl1(n41) );
	mux4_1 U122 ( .x(n285), .d0(D5_17), .d1(D13_17), .d2(D21_17), .d3(D29_17),
		.sl0(n8), .sl1(n37) );
	mux4_1 U123 ( .x(n317), .d0(D3_17), .d1(D11_17), .d2(D19_17), .d3(D27_17),
		.sl0(n8), .sl1(n39) );
	mux4_1 U124 ( .x(n253), .d0(D1_17), .d1(D9_17), .d2(D17_17), .d3(D25_17),
		.sl0(n16), .sl1(n35) );
	mux4_1 U125 ( .x(n189), .d0(D6_17), .d1(D14_17), .d2(D22_17), .d3(D30_17),
		.sl0(n15), .sl1(n33) );
	mux4_1 U126 ( .x(n125), .d0(D4_17), .d1(D12_17), .d2(D20_17), .d3(D28_17),
		.sl0(n14), .sl1(n29) );
	mux4_1 U127 ( .x(n157), .d0(D2_17), .d1(D10_17), .d2(D18_17), .d3(D26_17),
		.sl0(n11), .sl1(n31) );
	mux4_1 U128 ( .x(n93), .d0(D0_17), .d1(D8_17), .d2(D16_17), .d3(D24_17),
		.sl0(n13), .sl1(n27) );
	mux4_1 U129 ( .x(n358), .d0(D7_26), .d1(D15_26), .d2(D23_26), .d3(D31_26),
		.sl0(n7), .sl1(n41) );
	mux4_1 U13 ( .x(n203), .d0(D6_31), .d1(D14_31), .d2(D22_31), .d3(D30_31),
		.sl0(n16), .sl1(n33) );
	mux4_1 U130 ( .x(n294), .d0(D5_26), .d1(D13_26), .d2(D21_26), .d3(D29_26),
		.sl0(n8), .sl1(n37) );
	mux4_1 U131 ( .x(n326), .d0(D3_26), .d1(D11_26), .d2(D19_26), .d3(D27_26),
		.sl0(n18), .sl1(n39) );
	mux4_1 U132 ( .x(n262), .d0(D1_26), .d1(D9_26), .d2(D17_26), .d3(D25_26),
		.sl0(n16), .sl1(n35) );
	mux4_1 U133 ( .x(n198), .d0(D6_26), .d1(D14_26), .d2(D22_26), .d3(D30_26),
		.sl0(n10), .sl1(n33) );
	mux4_1 U134 ( .x(n134), .d0(D4_26), .d1(D12_26), .d2(D20_26), .d3(D28_26),
		.sl0(n14), .sl1(n29) );
	mux4_1 U135 ( .x(n166), .d0(D2_26), .d1(D10_26), .d2(D18_26), .d3(D26_26),
		.sl0(n21), .sl1(n31) );
	mux4_1 U136 ( .x(n102), .d0(D0_26), .d1(D8_26), .d2(D16_26), .d3(D24_26),
		.sl0(n13), .sl1(n27) );
	mux4_1 U137 ( .x(n340), .d0(D7_8), .d1(D15_8), .d2(D23_8), .d3(D31_8),
		.sl0(n24), .sl1(n40) );
	mux4_1 U138 ( .x(n276), .d0(D5_8), .d1(D13_8), .d2(D21_8), .d3(D29_8),
		.sl0(n23), .sl1(n36) );
	mux4_1 U139 ( .x(n308), .d0(D3_8), .d1(D11_8), .d2(D19_8), .d3(D27_8),
		.sl0(n8), .sl1(n38) );
	mux4_1 U14 ( .x(n139), .d0(D4_31), .d1(D12_31), .d2(D20_31), .d3(D28_31),
		.sl0(n14), .sl1(n29) );
	mux4_1 U140 ( .x(n244), .d0(D1_8), .d1(D9_8), .d2(D17_8), .d3(D25_8), .sl0(n16),
		.sl1(n34) );
	mux4_1 U141 ( .x(n180), .d0(D6_8), .d1(D14_8), .d2(D22_8), .d3(D30_8),
		.sl0(n21), .sl1(n32) );
	mux4_1 U142 ( .x(n116), .d0(D4_8), .d1(D12_8), .d2(D20_8), .d3(D28_8),
		.sl0(n20), .sl1(n28) );
	mux4_1 U143 ( .x(n148), .d0(D2_8), .d1(D10_8), .d2(D18_8), .d3(D26_8),
		.sl0(n11), .sl1(n30) );
	mux4_1 U144 ( .x(n84), .d0(D0_8), .d1(D8_8), .d2(D16_8), .d3(D24_8), .sl0(n19),
		.sl1(n26) );
	mux4_1 U145 ( .x(n339), .d0(D7_7), .d1(D15_7), .d2(D23_7), .d3(D31_7),
		.sl0(n18), .sl1(n40) );
	mux4_1 U146 ( .x(n275), .d0(D5_7), .d1(D13_7), .d2(D21_7), .d3(D29_7),
		.sl0(n16), .sl1(n36) );
	mux4_1 U147 ( .x(n307), .d0(D3_7), .d1(D11_7), .d2(D19_7), .d3(D27_7),
		.sl0(n17), .sl1(n38) );
	mux4_1 U148 ( .x(n243), .d0(D1_7), .d1(D9_7), .d2(D17_7), .d3(D25_7), .sl0(n16),
		.sl1(n34) );
	mux4_1 U149 ( .x(n179), .d0(D6_7), .d1(D14_7), .d2(D22_7), .d3(D30_7),
		.sl0(n15), .sl1(n32) );
	mux4_1 U15 ( .x(n171), .d0(D2_31), .d1(D10_31), .d2(D18_31), .d3(D26_31),
		.sl0(n15), .sl1(n31) );
	mux4_1 U150 ( .x(n115), .d0(D4_7), .d1(D12_7), .d2(D20_7), .d3(D28_7),
		.sl0(n14), .sl1(n28) );
	mux4_1 U151 ( .x(n147), .d0(D2_7), .d1(D10_7), .d2(D18_7), .d3(D26_7),
		.sl0(n20), .sl1(n30) );
	mux4_1 U152 ( .x(n83), .d0(D0_7), .d1(D8_7), .d2(D16_7), .d3(D24_7), .sl0(n12),
		.sl1(n26) );
	mux4_1 U153 ( .x(n362), .d0(D7_30), .d1(D15_30), .d2(D23_30), .d3(D31_30),
		.sl0(n19), .sl1(n41) );
	mux4_1 U154 ( .x(n298), .d0(D5_30), .d1(D13_30), .d2(D21_30), .d3(D29_30),
		.sl0(n23), .sl1(n37) );
	mux4_1 U155 ( .x(n330), .d0(D3_30), .d1(D11_30), .d2(D19_30), .d3(D27_30),
		.sl0(n7), .sl1(n39) );
	mux4_1 U156 ( .x(n266), .d0(D1_30), .d1(D9_30), .d2(D17_30), .d3(D25_30),
		.sl0(n16), .sl1(n35) );
	buf_3 U157 ( .x(n3), .a(S1) );
	mux4_1 U158 ( .x(n202), .d0(D6_30), .d1(D14_30), .d2(D22_30), .d3(D30_30),
		.sl0(n22), .sl1(n33) );
	mux4_1 U159 ( .x(n138), .d0(D4_30), .d1(D12_30), .d2(D20_30), .d3(D28_30),
		.sl0(n11), .sl1(n29) );
	mux4_1 U16 ( .x(n107), .d0(D0_31), .d1(D8_31), .d2(D16_31), .d3(D24_31),
		.sl0(n12), .sl1(n27) );
	mux4_1 U160 ( .x(n170), .d0(D2_30), .d1(D10_30), .d2(D18_30), .d3(D26_30),
		.sl0(n10), .sl1(n31) );
	mux4_1 U161 ( .x(n106), .d0(D0_30), .d1(D8_30), .d2(D16_30), .d3(D24_30),
		.sl0(n19), .sl1(n27) );
	mux4_2 U162 ( .x(n74), .d0(n106), .d1(n170), .d2(n138), .d3(n202), .sl0(n3),
		.sl1(n5) );
	mux4_1 U163 ( .x(n353), .d0(D7_21), .d1(D15_21), .d2(D23_21), .d3(D31_21),
		.sl0(n25), .sl1(n41) );
	mux4_1 U164 ( .x(n289), .d0(D5_21), .d1(D13_21), .d2(D21_21), .d3(D29_21),
		.sl0(n8), .sl1(n37) );
	mux4_1 U165 ( .x(n321), .d0(D3_21), .d1(D11_21), .d2(D19_21), .d3(D27_21),
		.sl0(n18), .sl1(n39) );
	mux4_1 U166 ( .x(n257), .d0(D1_21), .d1(D9_21), .d2(D17_21), .d3(D25_21),
		.sl0(n22), .sl1(n35) );
	mux4_1 U167 ( .x(n193), .d0(D6_21), .d1(D14_21), .d2(D22_21), .d3(D30_21),
		.sl0(n10), .sl1(n33) );
	mux4_1 U168 ( .x(n129), .d0(D4_21), .d1(D12_21), .d2(D20_21), .d3(D28_21),
		.sl0(n20), .sl1(n29) );
	mux4_1 U169 ( .x(n161), .d0(D2_21), .d1(D10_21), .d2(D18_21), .d3(D26_21),
		.sl0(n21), .sl1(n31) );
	mux4_1 U17 ( .x(n352), .d0(D7_20), .d1(D15_20), .d2(D23_20), .d3(D31_20),
		.sl0(n18), .sl1(n41) );
	mux4_1 U170 ( .x(n97), .d0(D0_21), .d1(D8_21), .d2(D16_21), .d3(D24_21),
		.sl0(n19), .sl1(n27) );
	mux4_1 U171 ( .x(n347), .d0(D7_15), .d1(D15_15), .d2(D23_15), .d3(D31_15),
		.sl0(n24), .sl1(n40) );
	mux4_1 U172 ( .x(n283), .d0(D5_15), .d1(D13_15), .d2(D21_15), .d3(D29_15),
		.sl0(n23), .sl1(n36) );
	mux4_1 U173 ( .x(n315), .d0(D3_15), .d1(D11_15), .d2(D19_15), .d3(D27_15),
		.sl0(n24), .sl1(n38) );
	mux4_1 U174 ( .x(n251), .d0(D1_15), .d1(D9_15), .d2(D17_15), .d3(D25_15),
		.sl0(n22), .sl1(n34) );
	mux4_1 U175 ( .x(n187), .d0(D6_15), .d1(D14_15), .d2(D22_15), .d3(D30_15),
		.sl0(n15), .sl1(n32) );
	mux4_1 U176 ( .x(n123), .d0(D4_15), .d1(D12_15), .d2(D20_15), .d3(D28_15),
		.sl0(n20), .sl1(n28) );
	mux4_1 U177 ( .x(n155), .d0(D2_15), .d1(D10_15), .d2(D18_15), .d3(D26_15),
		.sl0(n15), .sl1(n30) );
	mux4_1 U178 ( .x(n91), .d0(D0_15), .d1(D8_15), .d2(D16_15), .d3(D24_15),
		.sl0(n13), .sl1(n26) );
	mux4_1 U179 ( .x(n346), .d0(D7_14), .d1(D15_14), .d2(D23_14), .d3(D31_14),
		.sl0(n7), .sl1(n40) );
	mux4_1 U18 ( .x(n288), .d0(D5_20), .d1(D13_20), .d2(D21_20), .d3(D29_20),
		.sl0(n17), .sl1(n37) );
	mux4_1 U180 ( .x(n282), .d0(D5_14), .d1(D13_14), .d2(D21_14), .d3(D29_14),
		.sl0(n17), .sl1(n36) );
	mux4_1 U181 ( .x(n314), .d0(D3_14), .d1(D11_14), .d2(D19_14), .d3(D27_14),
		.sl0(n17), .sl1(n38) );
	mux4_1 U182 ( .x(n250), .d0(D1_14), .d1(D9_14), .d2(D17_14), .d3(D25_14),
		.sl0(n9), .sl1(n34) );
	mux4_2 U183 ( .x(n218), .d0(n250), .d1(n314), .d2(n282), .d3(n346), .sl0(n4),
		.sl1(n5) );
	mux4_1 U184 ( .x(n186), .d0(D6_14), .d1(D14_14), .d2(D22_14), .d3(D30_14),
		.sl0(n15), .sl1(n32) );
	mux4_1 U185 ( .x(n122), .d0(D4_14), .d1(D12_14), .d2(D20_14), .d3(D28_14),
		.sl0(n14), .sl1(n28) );
	mux4_1 U186 ( .x(n154), .d0(D2_14), .d1(D10_14), .d2(D18_14), .d3(D26_14),
		.sl0(n11), .sl1(n30) );
	mux4_1 U187 ( .x(n90), .d0(D0_14), .d1(D8_14), .d2(D16_14), .d3(D24_14),
		.sl0(n12), .sl1(n26) );
	mux4_2 U188 ( .x(n58), .d0(n90), .d1(n154), .d2(n122), .d3(n186), .sl0(n4),
		.sl1(n5) );
	mux4_1 U189 ( .x(n355), .d0(D7_23), .d1(D15_23), .d2(D23_23), .d3(D31_23),
		.sl0(n18), .sl1(n41) );
	mux4_1 U19 ( .x(n320), .d0(D3_20), .d1(D11_20), .d2(D19_20), .d3(D27_20),
		.sl0(n8), .sl1(n39) );
	mux4_1 U190 ( .x(n291), .d0(D5_23), .d1(D13_23), .d2(D21_23), .d3(D29_23),
		.sl0(n17), .sl1(n37) );
	mux4_1 U191 ( .x(n323), .d0(D3_23), .d1(D11_23), .d2(D19_23), .d3(D27_23),
		.sl0(n7), .sl1(n39) );
	mux4_1 U192 ( .x(n259), .d0(D1_23), .d1(D9_23), .d2(D17_23), .d3(D25_23),
		.sl0(n22), .sl1(n35) );
	mux4_1 U193 ( .x(n195), .d0(D6_23), .d1(D14_23), .d2(D22_23), .d3(D30_23),
		.sl0(n21), .sl1(n33) );
	mux4_1 U194 ( .x(n131), .d0(D4_23), .d1(D12_23), .d2(D20_23), .d3(D28_23),
		.sl0(n14), .sl1(n29) );
	mux4_1 U195 ( .x(n163), .d0(D2_23), .d1(D10_23), .d2(D18_23), .d3(D26_23),
		.sl0(n15), .sl1(n31) );
	mux4_1 U196 ( .x(n99), .d0(D0_23), .d1(D8_23), .d2(D16_23), .d3(D24_23),
		.sl0(n19), .sl1(n27) );
	mux4_1 U197 ( .x(n337), .d0(D7_5), .d1(D15_5), .d2(D23_5), .d3(D31_5),
		.sl0(n7), .sl1(n40) );
	mux4_1 U198 ( .x(n273), .d0(D5_5), .d1(D13_5), .d2(D21_5), .d3(D29_5),
		.sl0(n23), .sl1(n36) );
	mux4_1 U199 ( .x(n305), .d0(D3_5), .d1(D11_5), .d2(D19_5), .d3(D27_5),
		.sl0(n8), .sl1(n38) );
	mux4_1 U2 ( .x(n278), .d0(D5_10), .d1(D13_10), .d2(D21_10), .d3(D29_10),
		.sl0(n17), .sl1(n36) );
	mux4_1 U20 ( .x(n256), .d0(D1_20), .d1(D9_20), .d2(D17_20), .d3(D25_20),
		.sl0(n16), .sl1(n35) );
	mux4_1 U200 ( .x(n241), .d0(D1_5), .d1(D9_5), .d2(D17_5), .d3(D25_5), .sl0(n22),
		.sl1(n34) );
	mux4_1 U201 ( .x(n177), .d0(D6_5), .d1(D14_5), .d2(D22_5), .d3(D30_5),
		.sl0(n21), .sl1(n32) );
	mux4_1 U202 ( .x(n113), .d0(D4_5), .d1(D12_5), .d2(D20_5), .d3(D28_5),
		.sl0(n12), .sl1(n28) );
	mux4_1 U203 ( .x(n145), .d0(D2_5), .d1(D10_5), .d2(D18_5), .d3(D26_5),
		.sl0(n11), .sl1(n30) );
	mux4_1 U204 ( .x(n81), .d0(D0_5), .d1(D8_5), .d2(D16_5), .d3(D24_5), .sl0(n19),
		.sl1(n26) );
	mux4_1 U205 ( .x(n357), .d0(D7_25), .d1(D15_25), .d2(D23_25), .d3(D31_25),
		.sl0(n7), .sl1(n41) );
	mux4_1 U206 ( .x(n293), .d0(D5_25), .d1(D13_25), .d2(D21_25), .d3(D29_25),
		.sl0(n17), .sl1(n37) );
	mux4_1 U207 ( .x(n325), .d0(D3_25), .d1(D11_25), .d2(D19_25), .d3(D27_25),
		.sl0(n7), .sl1(n39) );
	mux4_1 U208 ( .x(n261), .d0(D1_25), .d1(D9_25), .d2(D17_25), .d3(D25_25),
		.sl0(n22), .sl1(n35) );
	mux4_1 U209 ( .x(n197), .d0(D6_25), .d1(D14_25), .d2(D22_25), .d3(D30_25),
		.sl0(n10), .sl1(n33) );
	mux4_1 U21 ( .x(n192), .d0(D6_20), .d1(D14_20), .d2(D22_20), .d3(D30_20),
		.sl0(n21), .sl1(n33) );
	mux4_1 U210 ( .x(n133), .d0(D4_25), .d1(D12_25), .d2(D20_25), .d3(D28_25),
		.sl0(n20), .sl1(n29) );
	mux4_1 U211 ( .x(n165), .d0(D2_25), .d1(D10_25), .d2(D18_25), .d3(D26_25),
		.sl0(n15), .sl1(n31) );
	mux4_1 U212 ( .x(n101), .d0(D0_25), .d1(D8_25), .d2(D16_25), .d3(D24_25),
		.sl0(n12), .sl1(n27) );
	mux4_1 U213 ( .x(n348), .d0(D7_16), .d1(D15_16), .d2(D23_16), .d3(D31_16),
		.sl0(n7), .sl1(n41) );
	mux4_1 U214 ( .x(n284), .d0(D5_16), .d1(D13_16), .d2(D21_16), .d3(D29_16),
		.sl0(n17), .sl1(n37) );
	mux4_1 U215 ( .x(n316), .d0(D3_16), .d1(D11_16), .d2(D19_16), .d3(D27_16),
		.sl0(n24), .sl1(n39) );
	mux4_1 U216 ( .x(n252), .d0(D1_16), .d1(D9_16), .d2(D17_16), .d3(D25_16),
		.sl0(n9), .sl1(n35) );
	mux4_1 U217 ( .x(n188), .d0(D6_16), .d1(D14_16), .d2(D22_16), .d3(D30_16),
		.sl0(n21), .sl1(n33) );
	mux4_1 U218 ( .x(n124), .d0(D4_16), .d1(D12_16), .d2(D20_16), .d3(D28_16),
		.sl0(n11), .sl1(n29) );
	mux4_1 U219 ( .x(n156), .d0(D2_16), .d1(D10_16), .d2(D18_16), .d3(D26_16),
		.sl0(n15), .sl1(n31) );
	mux4_1 U22 ( .x(n128), .d0(D4_20), .d1(D12_20), .d2(D20_20), .d3(D28_20),
		.sl0(n14), .sl1(n29) );
	mux4_1 U220 ( .x(n92), .d0(D0_16), .d1(D8_16), .d2(D16_16), .d3(D24_16),
		.sl0(n13), .sl1(n27) );
	mux4_1 U221 ( .x(n335), .d0(D7_3), .d1(D15_3), .d2(D23_3), .d3(D31_3),
		.sl0(n24), .sl1(n40) );
	mux4_1 U222 ( .x(n271), .d0(D5_3), .d1(D13_3), .d2(D21_3), .d3(D29_3),
		.sl0(n23), .sl1(n36) );
	mux4_1 U223 ( .x(n303), .d0(D3_3), .d1(D11_3), .d2(D19_3), .d3(D27_3),
		.sl0(n23), .sl1(n38) );
	mux4_1 U224 ( .x(n239), .d0(D1_3), .d1(D9_3), .d2(D17_3), .d3(D25_3), .sl0(n9),
		.sl1(n34) );
	mux4_1 U225 ( .x(n175), .d0(D6_3), .d1(D14_3), .d2(D22_3), .d3(D30_3),
		.sl0(n10), .sl1(n32) );
	mux4_1 U226 ( .x(n111), .d0(D4_3), .d1(D12_3), .d2(D20_3), .d3(D28_3),
		.sl0(n19), .sl1(n28) );
	mux4_1 U227 ( .x(n143), .d0(D2_3), .d1(D10_3), .d2(D18_3), .d3(D26_3),
		.sl0(n14), .sl1(n30) );
	mux4_1 U228 ( .x(n79), .d0(D0_3), .d1(D8_3), .d2(D16_3), .d3(D24_3), .sl0(n13),
		.sl1(n26) );
	buf_3 U229 ( .x(n25), .a(n43) );
	mux4_1 U23 ( .x(n160), .d0(D2_20), .d1(D10_20), .d2(D18_20), .d3(D26_20),
		.sl0(n11), .sl1(n31) );
	mux4_1 U230 ( .x(n360), .d0(D7_28), .d1(D15_28), .d2(D23_28), .d3(D31_28),
		.sl0(n25), .sl1(n41) );
	mux4_1 U231 ( .x(n296), .d0(D5_28), .d1(D13_28), .d2(D21_28), .d3(D29_28),
		.sl0(n17), .sl1(n37) );
	mux4_1 U232 ( .x(n328), .d0(D3_28), .d1(D11_28), .d2(D19_28), .d3(D27_28),
		.sl0(n24), .sl1(n39) );
	mux4_1 U233 ( .x(n264), .d0(D1_28), .d1(D9_28), .d2(D17_28), .d3(D25_28),
		.sl0(n9), .sl1(n35) );
	mux4_2 U234 ( .x(n232), .d0(n264), .d1(n328), .d2(n296), .d3(n360), .sl0(n3),
		.sl1(n5) );
	mux4_1 U235 ( .x(n200), .d0(D6_28), .d1(D14_28), .d2(D22_28), .d3(D30_28),
		.sl0(n16), .sl1(n33) );
	mux4_1 U236 ( .x(n136), .d0(D4_28), .d1(D12_28), .d2(D20_28), .d3(D28_28),
		.sl0(n20), .sl1(n29) );
	mux4_1 U237 ( .x(n168), .d0(D2_28), .d1(D10_28), .d2(D18_28), .d3(D26_28),
		.sl0(n21), .sl1(n31) );
	mux4_1 U238 ( .x(n104), .d0(D0_28), .d1(D8_28), .d2(D16_28), .d3(D24_28),
		.sl0(n13), .sl1(n27) );
	mux4_2 U239 ( .x(n72), .d0(n104), .d1(n168), .d2(n136), .d3(n200), .sl0(n3),
		.sl1(n5) );
	mux4_1 U24 ( .x(n96), .d0(D0_20), .d1(D8_20), .d2(D16_20), .d3(D24_20),
		.sl0(n12), .sl1(n27) );
	mux4_1 U240 ( .x(n361), .d0(D7_29), .d1(D15_29), .d2(D23_29), .d3(D31_29),
		.sl0(n25), .sl1(n41) );
	mux4_1 U241 ( .x(n297), .d0(D5_29), .d1(D13_29), .d2(D21_29), .d3(D29_29),
		.sl0(n23), .sl1(n37) );
	mux4_1 U242 ( .x(n329), .d0(D3_29), .d1(D11_29), .d2(D19_29), .d3(D27_29),
		.sl0(n24), .sl1(n39) );
	mux4_1 U243 ( .x(n265), .d0(D1_29), .d1(D9_29), .d2(D17_29), .d3(D25_29),
		.sl0(n22), .sl1(n35) );
	mux4_2 U244 ( .x(n233), .d0(n265), .d1(n329), .d2(n297), .d3(n361), .sl0(n3),
		.sl1(n5) );
	mux4_1 U245 ( .x(n201), .d0(D6_29), .d1(D14_29), .d2(D22_29), .d3(D30_29),
		.sl0(n22), .sl1(n33) );
	mux4_1 U246 ( .x(n137), .d0(D4_29), .d1(D12_29), .d2(D20_29), .d3(D28_29),
		.sl0(n11), .sl1(n29) );
	mux4_1 U247 ( .x(n169), .d0(D2_29), .d1(D10_29), .d2(D18_29), .d3(D26_29),
		.sl0(n10), .sl1(n31) );
	mux4_1 U248 ( .x(n105), .d0(D0_29), .d1(D8_29), .d2(D16_29), .d3(D24_29),
		.sl0(n19), .sl1(n27) );
	mux4_2 U249 ( .x(n73), .d0(n105), .d1(n169), .d2(n137), .d3(n201), .sl0(n3),
		.sl1(n5) );
	mux4_1 U25 ( .x(n343), .d0(D7_11), .d1(D15_11), .d2(D23_11), .d3(D31_11),
		.sl0(n7), .sl1(n40) );
	buf_3 U250 ( .x(n41), .a(S4) );
	buf_3 U251 ( .x(n37), .a(S4) );
	mux4_1 U252 ( .x(n295), .d0(D5_27), .d1(D13_27), .d2(D21_27), .d3(D29_27),
		.sl0(n23), .sl1(n37) );
	buf_3 U253 ( .x(n39), .a(S4) );
	buf_3 U254 ( .x(n35), .a(S4) );
	buf_3 U255 ( .x(n33), .a(S4) );
	buf_3 U256 ( .x(n29), .a(S4) );
	mux4_1 U257 ( .x(n135), .d0(D4_27), .d1(D12_27), .d2(D20_27), .d3(D28_27),
		.sl0(n11), .sl1(n29) );
	buf_3 U258 ( .x(n31), .a(S4) );
	mux4_1 U259 ( .x(n167), .d0(D2_27), .d1(D10_27), .d2(D18_27), .d3(D26_27),
		.sl0(n10), .sl1(n31) );
	mux4_1 U26 ( .x(n279), .d0(D5_11), .d1(D13_11), .d2(D21_11), .d3(D29_11),
		.sl0(n23), .sl1(n36) );
	buf_3 U260 ( .x(n27), .a(S4) );
	mux4_1 U261 ( .x(n103), .d0(D0_27), .d1(D8_27), .d2(D16_27), .d3(D24_27),
		.sl0(n13), .sl1(n27) );
	buf_3 U262 ( .x(n40), .a(S4) );
	mux4_1 U263 ( .x(n332), .d0(D7_0), .d1(D15_0), .d2(D23_0), .d3(D31_0),
		.sl0(n24), .sl1(n40) );
	buf_3 U264 ( .x(n36), .a(S4) );
	mux4_1 U265 ( .x(n268), .d0(D5_0), .d1(D13_0), .d2(D21_0), .d3(D29_0),
		.sl0(n16), .sl1(n36) );
	buf_3 U266 ( .x(n38), .a(S4) );
	mux4_1 U267 ( .x(n300), .d0(D3_0), .d1(D11_0), .d2(D19_0), .d3(D27_0),
		.sl0(n17), .sl1(n38) );
	buf_3 U268 ( .x(n34), .a(S4) );
	mux4_1 U269 ( .x(n236), .d0(D1_0), .d1(D9_0), .d2(D17_0), .d3(D25_0), .sl0(n16),
		.sl1(n34) );
	mux4_1 U27 ( .x(n311), .d0(D3_11), .d1(D11_11), .d2(D19_11), .d3(D27_11),
		.sl0(n8), .sl1(n38) );
	buf_3 U270 ( .x(n32), .a(S4) );
	mux4_1 U271 ( .x(n172), .d0(D6_0), .d1(D14_0), .d2(D22_0), .d3(D30_0),
		.sl0(n10), .sl1(n32) );
	buf_3 U272 ( .x(n28), .a(S4) );
	mux4_1 U273 ( .x(n108), .d0(D4_0), .d1(D12_0), .d2(D20_0), .d3(D28_0),
		.sl0(n12), .sl1(n28) );
	buf_3 U274 ( .x(n30), .a(S4) );
	mux4_1 U275 ( .x(n140), .d0(D2_0), .d1(D10_0), .d2(D18_0), .d3(D26_0),
		.sl0(n14), .sl1(n30) );
	buf_3 U276 ( .x(n26), .a(S4) );
	mux4_1 U277 ( .x(n76), .d0(D0_0), .d1(D8_0), .d2(D16_0), .d3(D24_0), .sl0(n13),
		.sl1(n26) );
	mux2_2 U278 ( .x(Z_10), .d0(n54), .sl(S0), .d1(n214) );
	mux2_2 U279 ( .x(Z_31), .d0(n75), .sl(S0), .d1(n235) );
	mux4_1 U28 ( .x(n247), .d0(D1_11), .d1(D9_11), .d2(D17_11), .d3(D25_11),
		.sl0(n16), .sl1(n34) );
	mux2_2 U280 ( .x(Z_20), .d0(n64), .sl(S0), .d1(n224) );
	mux2_2 U281 ( .x(Z_11), .d0(n55), .sl(S0), .d1(n215) );
	mux2_2 U282 ( .x(Z_1), .d0(n45), .sl(S0), .d1(n205) );
	mux2_2 U283 ( .x(Z_22), .d0(n66), .sl(S0), .d1(n226) );
	mux2_2 U284 ( .x(Z_6), .d0(n50), .sl(S0), .d1(n210) );
	mux2_2 U285 ( .x(Z_19), .d0(n63), .sl(S0), .d1(n223) );
	mux2_2 U286 ( .x(Z_9), .d0(n53), .sl(S0), .d1(n213) );
	mux2_2 U287 ( .x(Z_4), .d0(n48), .sl(S0), .d1(n208) );
	mux2_2 U288 ( .x(Z_24), .d0(n68), .sl(S0), .d1(n228) );
	mux2_2 U289 ( .x(Z_13), .d0(n57), .sl(S0), .d1(n217) );
	mux4_1 U29 ( .x(n183), .d0(D6_11), .d1(D14_11), .d2(D22_11), .d3(D30_11),
		.sl0(n21), .sl1(n32) );
	mux2_2 U290 ( .x(Z_18), .d0(n62), .sl(S0), .d1(n222) );
	mux2_2 U291 ( .x(Z_12), .d0(n56), .sl(S0), .d1(n216) );
	mux2_2 U292 ( .x(Z_17), .d0(n61), .sl(S0), .d1(n221) );
	mux2_2 U293 ( .x(Z_26), .d0(n70), .sl(S0), .d1(n230) );
	mux2_2 U294 ( .x(Z_8), .d0(n52), .sl(S0), .d1(n212) );
	mux2_2 U295 ( .x(Z_7), .d0(n51), .sl(S0), .d1(n211) );
	mux2_2 U296 ( .x(Z_30), .d0(n74), .sl(S0), .d1(n234) );
	mux2_2 U297 ( .x(Z_21), .d0(n65), .sl(S0), .d1(n225) );
	mux2_2 U298 ( .x(Z_15), .d0(n59), .sl(S0), .d1(n219) );
	mux2_2 U299 ( .x(Z_14), .d0(n58), .sl(S0), .d1(n218) );
	mux4_1 U3 ( .x(n310), .d0(D3_10), .d1(D11_10), .d2(D19_10), .d3(D27_10),
		.sl0(n24), .sl1(n38) );
	mux4_1 U30 ( .x(n119), .d0(D4_11), .d1(D12_11), .d2(D20_11), .d3(D28_11),
		.sl0(n12), .sl1(n28) );
	mux2_2 U300 ( .x(Z_23), .d0(n67), .sl(S0), .d1(n227) );
	mux2_2 U301 ( .x(Z_5), .d0(n49), .sl(S0), .d1(n209) );
	mux2_2 U302 ( .x(Z_25), .d0(n69), .sl(S0), .d1(n229) );
	mux2_2 U303 ( .x(Z_16), .d0(n60), .sl(S0), .d1(n220) );
	mux2_2 U304 ( .x(Z_3), .d0(n47), .sl(S0), .d1(n207) );
	mux2_2 U305 ( .x(Z_28), .d0(n72), .sl(S0), .d1(n232) );
	mux2_2 U306 ( .x(Z_29), .d0(n73), .sl(S0), .d1(n233) );
	mux2_2 U307 ( .x(Z_0), .d0(n44), .sl(S0), .d1(n204) );
	buf_10 U308 ( .x(n2), .a(S1) );
	buf_10 U309 ( .x(n1), .a(S1) );
	mux4_1 U31 ( .x(n151), .d0(D2_11), .d1(D10_11), .d2(D18_11), .d3(D26_11),
		.sl0(n20), .sl1(n30) );
	buf_4 U310 ( .x(n4), .a(S1) );
	buf_16 U313 ( .x(n7), .a(n43) );
	buf_16 U314 ( .x(n8), .a(n43) );
	buf_16 U315 ( .x(n9), .a(n43) );
	buf_16 U316 ( .x(n10), .a(n43) );
	buf_16 U317 ( .x(n11), .a(n43) );
	buf_16 U318 ( .x(n12), .a(n43) );
	buf_16 U319 ( .x(n13), .a(n43) );
	mux4_1 U32 ( .x(n87), .d0(D0_11), .d1(D8_11), .d2(D16_11), .d3(D24_11),
		.sl0(n12), .sl1(n26) );
	buf_16 U320 ( .x(n14), .a(n43) );
	buf_16 U321 ( .x(n15), .a(n43) );
	buf_16 U322 ( .x(n16), .a(n43) );
	buf_16 U323 ( .x(n17), .a(n43) );
	buf_16 U324 ( .x(n18), .a(n43) );
	buf_16 U325 ( .x(n19), .a(n43) );
	buf_16 U326 ( .x(n20), .a(n43) );
	buf_16 U327 ( .x(n21), .a(n43) );
	buf_16 U328 ( .x(n22), .a(n43) );
	buf_16 U329 ( .x(n23), .a(n43) );
	mux4_1 U33 ( .x(n333), .d0(D7_1), .d1(D15_1), .d2(D23_1), .d3(D31_1), .sl0(n18),
		.sl1(n40) );
	buf_16 U330 ( .x(n24), .a(n43) );
	inv_16 U331 ( .x(n43), .a(n42) );
	inv_16 U332 ( .x(n42), .a(S3) );
	mux2_4 U333 ( .x(Z_2), .d0(n46), .sl(S0), .d1(n206) );
	mux2_4 U334 ( .x(Z_27), .d0(n71), .sl(S0), .d1(n231) );
	mux4_3 U335 ( .x(n44), .d0(n76), .d1(n140), .d2(n108), .d3(n172), .sl0(n1),
		.sl1(n5) );
	mux4_3 U336 ( .x(n45), .d0(n77), .d1(n141), .d2(n109), .d3(n173), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U337 ( .x(n46), .d0(n78), .d1(n142), .d2(n110), .d3(n174), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U338 ( .x(n47), .d0(n79), .d1(n143), .d2(n111), .d3(n175), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U339 ( .x(n48), .d0(n80), .d1(n144), .d2(n112), .d3(n176), .sl0(n1),
		.sl1(n1425) );
	mux4_1 U34 ( .x(n269), .d0(D5_1), .d1(D13_1), .d2(D21_1), .d3(D29_1), .sl0(n9),
		.sl1(n36) );
	mux4_3 U340 ( .x(n49), .d0(n81), .d1(n145), .d2(n113), .d3(n177), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U341 ( .x(n50), .d0(n82), .d1(n146), .d2(n114), .d3(n178), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U342 ( .x(n51), .d0(n83), .d1(n147), .d2(n115), .d3(n179), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U343 ( .x(n52), .d0(n84), .d1(n148), .d2(n116), .d3(n180), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U344 ( .x(n53), .d0(n85), .d1(n149), .d2(n117), .d3(n181), .sl0(n3),
		.sl1(n1425) );
	mux4_3 U345 ( .x(n54), .d0(n86), .d1(n150), .d2(n118), .d3(n182), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U346 ( .x(n55), .d0(n87), .d1(n151), .d2(n119), .d3(n183), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U347 ( .x(n56), .d0(n88), .d1(n152), .d2(n120), .d3(n184), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U348 ( .x(n57), .d0(n89), .d1(n153), .d2(n121), .d3(n185), .sl0(n4),
		.sl1(n5) );
	mux4_3 U349 ( .x(n59), .d0(n91), .d1(n155), .d2(n123), .d3(n187), .sl0(n1),
		.sl1(n1425) );
	mux4_1 U35 ( .x(n301), .d0(D3_1), .d1(D11_1), .d2(D19_1), .d3(D27_1), .sl0(n17),
		.sl1(n38) );
	mux4_3 U350 ( .x(n60), .d0(n92), .d1(n156), .d2(n124), .d3(n188), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U351 ( .x(n61), .d0(n93), .d1(n157), .d2(n125), .d3(n189), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U352 ( .x(n62), .d0(n94), .d1(n158), .d2(n126), .d3(n190), .sl0(n4),
		.sl1(n5) );
	mux4_3 U353 ( .x(n63), .d0(n95), .d1(n159), .d2(n127), .d3(n191), .sl0(n3),
		.sl1(n1425) );
	mux4_3 U354 ( .x(n64), .d0(n96), .d1(n160), .d2(n128), .d3(n192), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U355 ( .x(n65), .d0(n97), .d1(n161), .d2(n129), .d3(n193), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U356 ( .x(n66), .d0(n98), .d1(n162), .d2(n130), .d3(n194), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U357 ( .x(n67), .d0(n99), .d1(n163), .d2(n131), .d3(n195), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U358 ( .x(n68), .d0(n100), .d1(n164), .d2(n132), .d3(n196), .sl0(n4),
		.sl1(n5) );
	mux4_3 U359 ( .x(n69), .d0(n101), .d1(n165), .d2(n133), .d3(n197), .sl0(n2),
		.sl1(n5) );
	mux4_1 U36 ( .x(n237), .d0(D1_1), .d1(D9_1), .d2(D17_1), .d3(D25_1), .sl0(n9),
		.sl1(n34) );
	mux4_3 U360 ( .x(n70), .d0(n102), .d1(n166), .d2(n134), .d3(n198), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U361 ( .x(n71), .d0(n103), .d1(n167), .d2(n135), .d3(n199), .sl0(n3),
		.sl1(n5) );
	mux4_3 U362 ( .x(n75), .d0(n107), .d1(n171), .d2(n139), .d3(n203), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U363 ( .x(n199), .d0(D6_27), .d1(D14_27), .d2(D22_27), .d3(D30_27),
		.sl0(n21), .sl1(n33) );
	mux4_3 U364 ( .x(n204), .d0(n236), .d1(n300), .d2(n268), .d3(n332), .sl0(n4),
		.sl1(n5) );
	mux4_3 U365 ( .x(n205), .d0(n237), .d1(n301), .d2(n269), .d3(n333), .sl0(n3),
		.sl1(n5) );
	mux4_3 U366 ( .x(n206), .d0(n238), .d1(n302), .d2(n270), .d3(n334), .sl0(n3),
		.sl1(n5) );
	mux4_3 U367 ( .x(n207), .d0(n239), .d1(n303), .d2(n271), .d3(n335), .sl0(n1),
		.sl1(n5) );
	mux4_3 U368 ( .x(n208), .d0(n240), .d1(n304), .d2(n272), .d3(n336), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U369 ( .x(n209), .d0(n241), .d1(n305), .d2(n273), .d3(n337), .sl0(n2),
		.sl1(n5) );
	mux4_1 U37 ( .x(n173), .d0(D6_1), .d1(D14_1), .d2(D22_1), .d3(D30_1), .sl0(n21),
		.sl1(n32) );
	mux4_3 U370 ( .x(n210), .d0(n242), .d1(n306), .d2(n274), .d3(n338), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U371 ( .x(n211), .d0(n243), .d1(n307), .d2(n275), .d3(n339), .sl0(n4),
		.sl1(n5) );
	mux4_3 U372 ( .x(n212), .d0(n244), .d1(n308), .d2(n276), .d3(n340), .sl0(n2),
		.sl1(n5) );
	mux4_3 U373 ( .x(n213), .d0(n245), .d1(n309), .d2(n277), .d3(n341), .sl0(n3),
		.sl1(n1425) );
	mux4_3 U374 ( .x(n214), .d0(n246), .d1(n310), .d2(n278), .d3(n342), .sl0(n3),
		.sl1(n1425) );
	mux4_3 U375 ( .x(n215), .d0(n247), .d1(n311), .d2(n279), .d3(n343), .sl0(n2),
		.sl1(n1425) );
	mux4_3 U376 ( .x(n216), .d0(n248), .d1(n312), .d2(n280), .d3(n344), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U377 ( .x(n217), .d0(n249), .d1(n313), .d2(n281), .d3(n345), .sl0(n1),
		.sl1(n5) );
	mux4_3 U378 ( .x(n219), .d0(n251), .d1(n315), .d2(n283), .d3(n347), .sl0(n4),
		.sl1(n1425) );
	mux4_3 U379 ( .x(n220), .d0(n252), .d1(n316), .d2(n284), .d3(n348), .sl0(n2),
		.sl1(n5) );
	mux4_1 U38 ( .x(n109), .d0(D4_1), .d1(D12_1), .d2(D20_1), .d3(D28_1), .sl0(n13),
		.sl1(n28) );
	mux4_3 U380 ( .x(n221), .d0(n253), .d1(n317), .d2(n285), .d3(n349), .sl0(n2),
		.sl1(n5) );
	mux4_3 U381 ( .x(n222), .d0(n254), .d1(n318), .d2(n286), .d3(n350), .sl0(n4),
		.sl1(n5) );
	mux4_3 U382 ( .x(n223), .d0(n255), .d1(n319), .d2(n287), .d3(n351), .sl0(n3),
		.sl1(n1425) );
	mux4_3 U383 ( .x(n224), .d0(n256), .d1(n320), .d2(n288), .d3(n352), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U384 ( .x(n225), .d0(n257), .d1(n321), .d2(n289), .d3(n353), .sl0(n1),
		.sl1(n5) );
	mux4_3 U385 ( .x(n226), .d0(n258), .d1(n322), .d2(n290), .d3(n354), .sl0(n4),
		.sl1(n5) );
	mux4_3 U386 ( .x(n227), .d0(n259), .d1(n323), .d2(n291), .d3(n355), .sl0(n1),
		.sl1(n5) );
	mux4_3 U387 ( .x(n228), .d0(n260), .d1(n324), .d2(n292), .d3(n356), .sl0(n1),
		.sl1(n5) );
	mux4_3 U388 ( .x(n229), .d0(n261), .d1(n325), .d2(n293), .d3(n357), .sl0(n1),
		.sl1(n5) );
	mux4_3 U389 ( .x(n230), .d0(n262), .d1(n326), .d2(n294), .d3(n358), .sl0(n4),
		.sl1(n5) );
	mux4_1 U39 ( .x(n141), .d0(D2_1), .d1(D10_1), .d2(D18_1), .d3(D26_1), .sl0(n20),
		.sl1(n30) );
	mux4_3 U390 ( .x(n231), .d0(n263), .d1(n327), .d2(n295), .d3(n359), .sl0(n3),
		.sl1(n5) );
	mux4_3 U391 ( .x(n234), .d0(n266), .d1(n330), .d2(n298), .d3(n362), .sl0(n3),
		.sl1(n5) );
	mux4_3 U392 ( .x(n235), .d0(n267), .d1(n331), .d2(n299), .d3(n363), .sl0(n1),
		.sl1(n1425) );
	mux4_3 U393 ( .x(n263), .d0(D1_27), .d1(D9_27), .d2(D17_27), .d3(D25_27),
		.sl0(n22), .sl1(n35) );
	mux4_3 U394 ( .x(n327), .d0(D3_27), .d1(D11_27), .d2(D19_27), .d3(D27_27),
		.sl0(n7), .sl1(n39) );
	mux4_3 U395 ( .x(n359), .d0(D7_27), .d1(D15_27), .d2(D23_27), .d3(D31_27),
		.sl0(n19), .sl1(n41) );
	buf_3 U396 ( .x(n1425), .a(S2) );
	buf_3 U397 ( .x(n5), .a(S2) );
	mux4_1 U4 ( .x(n246), .d0(D1_10), .d1(D9_10), .d2(D17_10), .d3(D25_10),
		.sl0(n9), .sl1(n34) );
	mux4_1 U40 ( .x(n77), .d0(D0_1), .d1(D8_1), .d2(D16_1), .d3(D24_1), .sl0(n13),
		.sl1(n26) );
	mux4_1 U41 ( .x(n354), .d0(D7_22), .d1(D15_22), .d2(D23_22), .d3(D31_22),
		.sl0(n7), .sl1(n41) );
	mux4_1 U42 ( .x(n290), .d0(D5_22), .d1(D13_22), .d2(D21_22), .d3(D29_22),
		.sl0(n23), .sl1(n37) );
	mux4_1 U43 ( .x(n322), .d0(D3_22), .d1(D11_22), .d2(D19_22), .d3(D27_22),
		.sl0(n24), .sl1(n39) );
	mux4_1 U44 ( .x(n258), .d0(D1_22), .d1(D9_22), .d2(D17_22), .d3(D25_22),
		.sl0(n9), .sl1(n35) );
	mux4_1 U45 ( .x(n194), .d0(D6_22), .d1(D14_22), .d2(D22_22), .d3(D30_22),
		.sl0(n10), .sl1(n33) );
	mux4_1 U46 ( .x(n130), .d0(D4_22), .d1(D12_22), .d2(D20_22), .d3(D28_22),
		.sl0(n11), .sl1(n29) );
	mux4_1 U47 ( .x(n162), .d0(D2_22), .d1(D10_22), .d2(D18_22), .d3(D26_22),
		.sl0(n10), .sl1(n31) );
	mux4_1 U48 ( .x(n98), .d0(D0_22), .d1(D8_22), .d2(D16_22), .d3(D24_22),
		.sl0(n13), .sl1(n27) );
	mux4_1 U49 ( .x(n334), .d0(D7_2), .d1(D15_2), .d2(D23_2), .d3(D31_2), .sl0(n24),
		.sl1(n40) );
	mux4_1 U5 ( .x(n182), .d0(D6_10), .d1(D14_10), .d2(D22_10), .d3(D30_10),
		.sl0(n15), .sl1(n32) );
	mux4_1 U50 ( .x(n270), .d0(D5_2), .d1(D13_2), .d2(D21_2), .d3(D29_2), .sl0(n22),
		.sl1(n36) );
	mux4_1 U51 ( .x(n302), .d0(D3_2), .d1(D11_2), .d2(D19_2), .d3(D27_2), .sl0(n17),
		.sl1(n38) );
	mux4_1 U52 ( .x(n238), .d0(D1_2), .d1(D9_2), .d2(D17_2), .d3(D25_2), .sl0(n22),
		.sl1(n34) );
	mux4_1 U53 ( .x(n174), .d0(D6_2), .d1(D14_2), .d2(D22_2), .d3(D30_2), .sl0(n10),
		.sl1(n32) );
	mux4_1 U54 ( .x(n110), .d0(D4_2), .d1(D12_2), .d2(D20_2), .d3(D28_2), .sl0(n12),
		.sl1(n28) );
	mux4_1 U55 ( .x(n142), .d0(D2_2), .d1(D10_2), .d2(D18_2), .d3(D26_2), .sl0(n11),
		.sl1(n30) );
	mux4_1 U56 ( .x(n78), .d0(D0_2), .d1(D8_2), .d2(D16_2), .d3(D24_2), .sl0(n12),
		.sl1(n26) );
	mux4_1 U57 ( .x(n338), .d0(D7_6), .d1(D15_6), .d2(D23_6), .d3(D31_6), .sl0(n18),
		.sl1(n40) );
	mux4_1 U58 ( .x(n274), .d0(D5_6), .d1(D13_6), .d2(D21_6), .d3(D29_6), .sl0(n9),
		.sl1(n36) );
	mux4_1 U59 ( .x(n306), .d0(D3_6), .d1(D11_6), .d2(D19_6), .d3(D27_6), .sl0(n23),
		.sl1(n38) );
	mux4_1 U6 ( .x(n118), .d0(D4_10), .d1(D12_10), .d2(D20_10), .d3(D28_10),
		.sl0(n14), .sl1(n28) );
	mux4_1 U60 ( .x(n242), .d0(D1_6), .d1(D9_6), .d2(D17_6), .d3(D25_6), .sl0(n16),
		.sl1(n34) );
	mux4_1 U61 ( .x(n178), .d0(D6_6), .d1(D14_6), .d2(D22_6), .d3(D30_6), .sl0(n10),
		.sl1(n32) );
	mux4_1 U62 ( .x(n114), .d0(D4_6), .d1(D12_6), .d2(D20_6), .d3(D28_6), .sl0(n19),
		.sl1(n28) );
	mux4_1 U63 ( .x(n146), .d0(D2_6), .d1(D10_6), .d2(D18_6), .d3(D26_6), .sl0(n14),
		.sl1(n30) );
	mux4_1 U64 ( .x(n82), .d0(D0_6), .d1(D8_6), .d2(D16_6), .d3(D24_6), .sl0(n12),
		.sl1(n26) );
	mux4_1 U65 ( .x(n351), .d0(D7_19), .d1(D15_19), .d2(D23_19), .d3(D31_19),
		.sl0(n7), .sl1(n41) );
	mux4_1 U66 ( .x(n287), .d0(D5_19), .d1(D13_19), .d2(D21_19), .d3(D29_19),
		.sl0(n17), .sl1(n37) );
	mux4_1 U67 ( .x(n319), .d0(D3_19), .d1(D11_19), .d2(D19_19), .d3(D27_19),
		.sl0(n24), .sl1(n39) );
	mux4_1 U68 ( .x(n255), .d0(D1_19), .d1(D9_19), .d2(D17_19), .d3(D25_19),
		.sl0(n9), .sl1(n35) );
	mux4_1 U69 ( .x(n191), .d0(D6_19), .d1(D14_19), .d2(D22_19), .d3(D30_19),
		.sl0(n10), .sl1(n33) );
	mux4_1 U7 ( .x(n150), .d0(D2_10), .d1(D10_10), .d2(D18_10), .d3(D26_10),
		.sl0(n14), .sl1(n30) );
	mux4_1 U70 ( .x(n127), .d0(D4_19), .d1(D12_19), .d2(D20_19), .d3(D28_19),
		.sl0(n11), .sl1(n29) );
	mux4_1 U71 ( .x(n159), .d0(D2_19), .d1(D10_19), .d2(D18_19), .d3(D26_19),
		.sl0(n21), .sl1(n31) );
	mux4_1 U72 ( .x(n95), .d0(D0_19), .d1(D8_19), .d2(D16_19), .d3(D24_19),
		.sl0(n12), .sl1(n27) );
	mux4_1 U73 ( .x(n341), .d0(D7_9), .d1(D15_9), .d2(D23_9), .d3(D31_9), .sl0(n24),
		.sl1(n40) );
	mux4_1 U74 ( .x(n277), .d0(D5_9), .d1(D13_9), .d2(D21_9), .d3(D29_9), .sl0(n8),
		.sl1(n36) );
	mux4_1 U75 ( .x(n309), .d0(D3_9), .d1(D11_9), .d2(D19_9), .d3(D27_9), .sl0(n23),
		.sl1(n38) );
	mux4_1 U76 ( .x(n245), .d0(D1_9), .d1(D9_9), .d2(D17_9), .d3(D25_9), .sl0(n22),
		.sl1(n34) );
	mux4_1 U77 ( .x(n181), .d0(D6_9), .d1(D14_9), .d2(D22_9), .d3(D30_9), .sl0(n10),
		.sl1(n32) );
	mux4_1 U78 ( .x(n117), .d0(D4_9), .d1(D12_9), .d2(D20_9), .d3(D28_9), .sl0(n20),
		.sl1(n28) );
	mux4_1 U79 ( .x(n149), .d0(D2_9), .d1(D10_9), .d2(D18_9), .d3(D26_9), .sl0(n14),
		.sl1(n30) );
	mux4_1 U8 ( .x(n86), .d0(D0_10), .d1(D8_10), .d2(D16_10), .d3(D24_10),
		.sl0(n19), .sl1(n26) );
	mux4_1 U80 ( .x(n85), .d0(D0_9), .d1(D8_9), .d2(D16_9), .d3(D24_9), .sl0(n13),
		.sl1(n26) );
	mux4_1 U81 ( .x(n336), .d0(D7_4), .d1(D15_4), .d2(D23_4), .d3(D31_4), .sl0(n7),
		.sl1(n40) );
	mux4_1 U82 ( .x(n272), .d0(D5_4), .d1(D13_4), .d2(D21_4), .d3(D29_4), .sl0(n9),
		.sl1(n36) );
	mux4_1 U83 ( .x(n304), .d0(D3_4), .d1(D11_4), .d2(D19_4), .d3(D27_4), .sl0(n8),
		.sl1(n38) );
	mux4_1 U84 ( .x(n240), .d0(D1_4), .d1(D9_4), .d2(D17_4), .d3(D25_4), .sl0(n9),
		.sl1(n34) );
	mux4_1 U85 ( .x(n176), .d0(D6_4), .d1(D14_4), .d2(D22_4), .d3(D30_4), .sl0(n15),
		.sl1(n32) );
	mux4_1 U86 ( .x(n112), .d0(D4_4), .d1(D12_4), .d2(D20_4), .d3(D28_4), .sl0(n13),
		.sl1(n28) );
	mux4_1 U87 ( .x(n144), .d0(D2_4), .d1(D10_4), .d2(D18_4), .d3(D26_4), .sl0(n20),
		.sl1(n30) );
	mux4_1 U88 ( .x(n80), .d0(D0_4), .d1(D8_4), .d2(D16_4), .d3(D24_4), .sl0(n19),
		.sl1(n26) );
	mux4_1 U89 ( .x(n356), .d0(D7_24), .d1(D15_24), .d2(D23_24), .d3(D31_24),
		.sl0(n18), .sl1(n41) );
	mux4_1 U9 ( .x(n363), .d0(D7_31), .d1(D15_31), .d2(D23_31), .d3(D31_31),
		.sl0(n25), .sl1(n41) );
	mux4_1 U90 ( .x(n292), .d0(D5_24), .d1(D13_24), .d2(D21_24), .d3(D29_24),
		.sl0(n23), .sl1(n37) );
	mux4_1 U91 ( .x(n324), .d0(D3_24), .d1(D11_24), .d2(D19_24), .d3(D27_24),
		.sl0(n18), .sl1(n39) );
	mux4_1 U92 ( .x(n260), .d0(D1_24), .d1(D9_24), .d2(D17_24), .d3(D25_24),
		.sl0(n9), .sl1(n35) );
	mux4_1 U93 ( .x(n196), .d0(D6_24), .d1(D14_24), .d2(D22_24), .d3(D30_24),
		.sl0(n21), .sl1(n33) );
	mux4_1 U94 ( .x(n132), .d0(D4_24), .d1(D12_24), .d2(D20_24), .d3(D28_24),
		.sl0(n14), .sl1(n29) );
	mux4_1 U95 ( .x(n164), .d0(D2_24), .d1(D10_24), .d2(D18_24), .d3(D26_24),
		.sl0(n15), .sl1(n31) );
	mux4_1 U96 ( .x(n100), .d0(D0_24), .d1(D8_24), .d2(D16_24), .d3(D24_24),
		.sl0(n12), .sl1(n27) );
	mux4_1 U97 ( .x(n345), .d0(D7_13), .d1(D15_13), .d2(D23_13), .d3(D31_13),
		.sl0(n18), .sl1(n40) );
	mux4_1 U98 ( .x(n281), .d0(D5_13), .d1(D13_13), .d2(D21_13), .d3(D29_13),
		.sl0(n8), .sl1(n36) );
	mux4_1 U99 ( .x(n313), .d0(D3_13), .d1(D11_13), .d2(D19_13), .d3(D27_13),
		.sl0(n17), .sl1(n38) );

endmodule


module ID_DW01_sub_32_2_test_1 (  A, B, CI, DIFF, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] DIFF;

wire A_0, A_1, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
	n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
	n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
	n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
	n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
	n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
	n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
	n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
	n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
	n206, n50, n52, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65,
	n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79,
	n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
	n94, n95, n96, n97, n98, n99;

	assign A_1 = A[1];
	assign A_0 = A[0];
	assign DIFF[1] = A_1;
	assign DIFF[0] = A_0;

	nor2_1 U10 ( .x(n176), .a(A[29]), .b(A[28]) );
	nor2i_2 U100 ( .x(n67), .a(n157), .b(n81) );
	nor2_1 U101 ( .x(n170), .a(A[9]), .b(A[8]) );
	nor2_1 U102 ( .x(n155), .a(A[6]), .b(A[10]) );
	oa21_4 U103 ( .x(DIFF[6]), .a(n63), .b(n130), .c(n62) );
	nand2_0 U104 ( .x(n62), .a(n129), .b(n71) );
	nand2_1 U105 ( .x(n63), .a(n167), .b(n64) );
	inv_1 U106 ( .x(n64), .a(n136) );
	oai21_5 U108 ( .x(DIFF[17]), .a(n95), .b(n96), .c(n97) );
	inv_0 U109 ( .x(n90), .a(A[15]) );
	nand2i_2 U11 ( .x(n177), .a(A[27]), .b(n124) );
	nand3i_1 U110 ( .x(n142), .a(A[15]), .b(n169), .c(n137) );
	mux2_2 U111 ( .x(n65), .d0(n161), .sl(n167), .d1(n136) );
	nand2i_1 U112 ( .x(n136), .a(A[4]), .b(n137) );
	inv_1 U113 ( .x(n161), .a(n70) );
	nand2i_0 U114 ( .x(n162), .a(A[8]), .b(n135) );
	inv_2 U115 ( .x(DIFF[2]), .a(A[2]) );
	nor2_0 U116 ( .x(n165), .a(A[2]), .b(A[3]) );
	inv_0 U118 ( .x(n104), .a(A[20]) );
	oai21_1 U119 ( .x(DIFF[4]), .a(n68), .b(n69), .c(n70) );
	inv_0 U120 ( .x(n129), .a(A[6]) );
	nand2i_2 U121 ( .x(n199), .a(A[12]), .b(n157) );
	inv_0 U122 ( .x(n87), .a(A[13]) );
	nand2i_2 U123 ( .x(n70), .a(A[4]), .b(n160) );
	nor2_1 U124 ( .x(n173), .a(A[10]), .b(A[13]) );
	nand3i_1 U125 ( .x(n174), .a(A[14]), .b(n99), .c(n173) );
	nor2_1 U126 ( .x(n188), .a(A[13]), .b(A[14]) );
	inv_2 U127 ( .x(n149), .a(A[3]) );
	nand2i_0 U129 ( .x(n198), .a(A[11]), .b(n197) );
	nand3i_0 U130 ( .x(n189), .a(A[11]), .b(n188), .c(n187) );
	nand4i_1 U131 ( .x(n182), .a(A[11]), .b(n181), .c(n180), .d(n179) );
	nor2_0 U133 ( .x(n193), .a(A[9]), .b(A[8]) );
	nand4i_1 U134 ( .x(n72), .a(A[7]), .b(n165), .c(n166), .d(n69) );
	nand2i_0 U135 ( .x(n164), .a(A[7]), .b(n163) );
	inv_0 U136 ( .x(n84), .a(A[12]) );
	nor2_0 U137 ( .x(n197), .a(A[12]), .b(A[13]) );
	nor2_0 U138 ( .x(n191), .a(A[12]), .b(A[11]) );
	nor2_0 U139 ( .x(n184), .a(A[12]), .b(A[11]) );
	nand2i_0 U14 ( .x(n83), .a(n157), .b(n81) );
	nor2_0 U140 ( .x(n180), .a(A[15]), .b(A[12]) );
	inv_0 U141 ( .x(n167), .a(A[5]) );
	nor2_0 U142 ( .x(n166), .a(A[6]), .b(A[5]) );
	nor3_0 U143 ( .x(n195), .a(A[4]), .b(A[6]), .c(A[5]) );
	oai21_4 U146 ( .x(DIFF[9]), .a(n76), .b(n77), .c(n78) );
	oai21_4 U147 ( .x(DIFF[13]), .a(n86), .b(n87), .c(n88) );
	oai21_4 U148 ( .x(DIFF[24]), .a(n112), .b(n113), .c(n114) );
	nand2i_4 U149 ( .x(n139), .a(n140), .b(n141) );
	nor2i_1 U15 ( .x(n192), .a(n191), .b(n190) );
	and3i_3 U150 ( .x(n144), .a(n174), .b(n172), .c(n171) );
	inv_5 U151 ( .x(n68), .a(n200) );
	nand2i_4 U152 ( .x(n74), .a(n162), .b(n130) );
	nand2i_4 U153 ( .x(n78), .a(n164), .b(n130) );
	nand2i_4 U154 ( .x(n85), .a(n199), .b(n201) );
	inv_5 U155 ( .x(n86), .a(n85) );
	nand2i_4 U156 ( .x(n88), .a(n198), .b(n201) );
	inv_5 U157 ( .x(n98), .a(n97) );
	nand2i_4 U158 ( .x(n101), .a(A[19]), .b(n146) );
	inv_5 U159 ( .x(n202), .a(n105) );
	nand2i_0 U16 ( .x(n194), .a(A[7]), .b(n193) );
	nand2_5 U160 ( .x(n106), .a(n202), .b(n153) );
	nand2_5 U161 ( .x(n110), .a(n203), .b(n151) );
	nand2i_4 U162 ( .x(n114), .a(n178), .b(n203) );
	nand2i_4 U165 ( .x(n122), .a(n150), .b(n120) );
	nand2i_4 U166 ( .x(n111), .a(n151), .b(n109) );
	nand2i_4 U167 ( .x(n107), .a(n153), .b(n105) );
	nand2_5 U168 ( .x(DIFF[19]), .a(n101), .b(n102) );
	oai21_5 U169 ( .x(DIFF[28]), .a(n123), .b(n124), .c(n125) );
	nand4i_1 U17 ( .x(n89), .a(n194), .b(n192), .c(n196), .d(n195) );
	oai21_5 U170 ( .x(DIFF[29]), .a(n126), .b(n127), .c(n128) );
	exnor2_5 U171 ( .x(DIFF[30]), .a(n159), .b(n132) );
	nand2_5 U172 ( .x(DIFF[8]), .a(n74), .b(n75) );
	nand2i_5 U173 ( .x(n91), .a(n189), .b(n201) );
	nand2i_5 U174 ( .x(n94), .a(n186), .b(n201) );
	nand2i_5 U175 ( .x(n97), .a(n182), .b(n201) );
	nand3i_5 U176 ( .x(n100), .a(n142), .b(n143), .c(n144) );
	nand2i_6 U178 ( .x(n105), .a(n152), .b(n146) );
	inv_2 U18 ( .x(n69), .a(A[4]) );
	inv_6 U180 ( .x(n123), .a(n121) );
	nand2i_6 U181 ( .x(n125), .a(n177), .b(n148) );
	nand2i_6 U182 ( .x(n128), .a(n147), .b(n148) );
	nor2i_5 U183 ( .x(n143), .a(n170), .b(n199) );
	nand2_3 U185 ( .x(n145), .a(n175), .b(n119) );
	nor2_1 U187 ( .x(n133), .a(A[5]), .b(A[6]) );
	ao21_4 U188 ( .x(DIFF[26]), .a(n117), .b(A[26]), .c(n148) );
	inv_2 U189 ( .x(n118), .a(n117) );
	inv_4 U190 ( .x(n119), .a(A[26]) );
	nand2i_4 U191 ( .x(n120), .a(n145), .b(n146) );
	inv_7 U192 ( .x(n148), .a(n120) );
	nand2i_1 U193 ( .x(n117), .a(n139), .b(n146) );
	nand3_1 U194 ( .x(n71), .a(n69), .b(n133), .c(n134) );
	nor2_0 U195 ( .x(n172), .a(A[5]), .b(A[6]) );
	nand2_1 U196 ( .x(n102), .a(A[19]), .b(n100) );
	inv_8 U197 ( .x(n146), .a(n100) );
	oai21_2 U198 ( .x(DIFF[20]), .a(n104), .b(n103), .c(n105) );
	nand4_5 U199 ( .x(n81), .a(n68), .b(n50), .c(n155), .d(n156) );
	nand2i_2 U20 ( .x(n75), .a(n66), .b(n72) );
	inv_4 U200 ( .x(n130), .a(n71) );
	nand2i_1 U201 ( .x(n73), .a(n135), .b(n71) );
	aoi21_6 U202 ( .x(n204), .a(n206), .b(n205), .c(n118) );
	inv_7 U203 ( .x(DIFF[25]), .a(n204) );
	inv_2 U204 ( .x(n205), .a(n116) );
	inv_10 U205 ( .x(n206), .a(n115) );
	inv_7 U206 ( .x(n115), .a(n114) );
	nor2_3 U207 ( .x(n56), .a(A[20]), .b(A[19]) );
	nand2i_2 U208 ( .x(n152), .a(A[20]), .b(n154) );
	nor2_2 U209 ( .x(n168), .a(A[25]), .b(A[24]) );
	inv_2 U21 ( .x(n175), .a(n139) );
	nand2i_0 U210 ( .x(n178), .a(A[24]), .b(n151) );
	inv_6 U211 ( .x(n96), .a(A[17]) );
	nor2_1 U212 ( .x(n179), .a(A[17]), .b(A[16]) );
	inv_3 U213 ( .x(n66), .a(A[8]) );
	nor2_1 U214 ( .x(n163), .a(A[9]), .b(A[8]) );
	inv_4 U215 ( .x(n108), .a(A[22]) );
	nand3_1 U22 ( .x(n186), .a(n185), .b(n183), .c(n184) );
	nor2_0 U24 ( .x(n181), .a(A[14]), .b(A[13]) );
	nor2i_1 U26 ( .x(n131), .a(n132), .b(n128) );
	inv_1 U27 ( .x(n80), .a(A[10]) );
	nand2_3 U28 ( .x(n121), .a(n148), .b(n150) );
	nand2_2 U29 ( .x(DIFF[27]), .a(n121), .b(n122) );
	nand2_2 U30 ( .x(DIFF[7]), .a(n72), .b(n73) );
	inv_2 U31 ( .x(n126), .a(n125) );
	inv_2 U34 ( .x(n95), .a(n94) );
	inv_2 U35 ( .x(n92), .a(n91) );
	oai21_1 U36 ( .x(DIFF[16]), .a(n92), .b(n93), .c(n94) );
	nand2_2 U37 ( .x(DIFF[11]), .a(n82), .b(n83) );
	inv_2 U38 ( .x(n82), .a(n67) );
	inv_5 U39 ( .x(n203), .a(n109) );
	nor2_0 U4 ( .x(n187), .a(A[15]), .b(A[12]) );
	oai21_3 U40 ( .x(DIFF[15]), .a(n57), .b(n90), .c(n91) );
	inv_2 U41 ( .x(n79), .a(n78) );
	inv_2 U42 ( .x(n76), .a(n74) );
	inv_2 U44 ( .x(n112), .a(n110) );
	nand2_2 U45 ( .x(DIFF[21]), .a(n106), .b(n107) );
	oai21_2 U46 ( .x(DIFF[18]), .a(n98), .b(n99), .c(n100) );
	nand2_2 U47 ( .x(DIFF[23]), .a(n110), .b(n111) );
	inv_2 U48 ( .x(n159), .a(n128) );
	exnor2_1 U49 ( .x(DIFF[31]), .a(n131), .b(n158) );
	nand2i_2 U5 ( .x(n190), .a(A[2]), .b(n149) );
	inv_3 U50 ( .x(DIFF[5]), .a(n65) );
	inv_2 U51 ( .x(n99), .a(A[18]) );
	inv_0 U52 ( .x(n113), .a(A[24]) );
	inv_0 U53 ( .x(n116), .a(A[25]) );
	inv_2 U54 ( .x(n151), .a(A[23]) );
	inv_2 U55 ( .x(n135), .a(A[7]) );
	inv_2 U57 ( .x(n150), .a(A[27]) );
	inv_2 U58 ( .x(n124), .a(A[28]) );
	inv_2 U59 ( .x(n127), .a(A[29]) );
	nand2i_2 U6 ( .x(n140), .a(A[23]), .b(n168) );
	inv_2 U60 ( .x(n132), .a(A[30]) );
	inv_2 U61 ( .x(n158), .a(A[31]) );
	and3_5 U62 ( .x(n50), .a(n135), .b(n66), .c(n77) );
	ao21_6 U63 ( .x(DIFF[22]), .a(n106), .b(n52), .c(n203) );
	inv_2 U64 ( .x(n52), .a(n108) );
	nand2i_4 U66 ( .x(n109), .a(n138), .b(n146) );
	oai21_3 U69 ( .x(DIFF[12]), .a(n84), .b(n67), .c(n85) );
	nor2_0 U7 ( .x(n185), .a(A[13]), .b(A[14]) );
	nor2_1 U70 ( .x(n156), .a(A[4]), .b(A[5]) );
	inv_3 U71 ( .x(n77), .a(A[9]) );
	inv_5 U72 ( .x(n57), .a(n89) );
	nand3_2 U73 ( .x(n138), .a(n153), .b(n108), .c(n56) );
	or2_2 U75 ( .x(n55), .a(A[7]), .b(A[4]) );
	inv_2 U76 ( .x(n171), .a(n55) );
	inv_10 U77 ( .x(n201), .a(n81) );
	inv_2 U8 ( .x(n141), .a(n138) );
	nor2_0 U81 ( .x(n183), .a(A[16]), .b(A[15]) );
	inv_0 U82 ( .x(n93), .a(A[16]) );
	nor2_3 U83 ( .x(n137), .a(A[2]), .b(A[3]) );
	nor2_1 U84 ( .x(n134), .a(A[2]), .b(A[3]) );
	inv_0 U85 ( .x(n154), .a(A[19]) );
	ao21_3 U86 ( .x(DIFF[14]), .a(n88), .b(A[14]), .c(n57) );
	nand2i_2 U87 ( .x(n58), .a(A[16]), .b(n96) );
	inv_2 U88 ( .x(n169), .a(n58) );
	oai21_1 U89 ( .x(DIFF[3]), .a(n149), .b(n59), .c(n200) );
	nand2i_2 U9 ( .x(n147), .a(A[27]), .b(n176) );
	inv_0 U90 ( .x(n59), .a(A[2]) );
	and3_2 U91 ( .x(n196), .a(n60), .b(n80), .c(n61) );
	inv_0 U92 ( .x(n60), .a(A[13]) );
	inv_0 U93 ( .x(n61), .a(A[14]) );
	inv_6 U94 ( .x(n103), .a(n101) );
	nand2i_4 U95 ( .x(n200), .a(A[2]), .b(n149) );
	nor2_1 U96 ( .x(n160), .a(A[2]), .b(A[3]) );
	inv_2 U97 ( .x(n153), .a(A[21]) );
	inv_5 U98 ( .x(n157), .a(A[11]) );
	oai21_1 U99 ( .x(DIFF[10]), .a(n79), .b(n80), .c(n81) );

endmodule


module ID_DW01_sub_32_0_test_1 (  A, B, CI, DIFF, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] DIFF;

wire A_0, A_1, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
	n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
	n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
	n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
	n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
	n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
	n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
	n182, n183, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61,
	n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n75, n76,
	n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
	n91, n92, n93, n94, n95, n96, n97, n98, n99;

	assign A_1 = A[1];
	assign A_0 = A[0];
	assign DIFF[1] = A_1;
	assign DIFF[0] = A_0;

	nand2i_1 U10 ( .x(n123), .a(n162), .b(n121) );
	nand2_4 U100 ( .x(n110), .a(n177), .b(n116) );
	nor2i_2 U101 ( .x(n130), .a(n131), .b(n132) );
	nand2i_2 U102 ( .x(n127), .a(n160), .b(n124) );
	nor2i_5 U103 ( .x(n57), .a(n162), .b(n121) );
	nand2i_2 U104 ( .x(n125), .a(n161), .b(n55) );
	nand2_5 U105 ( .x(DIFF[25]), .a(n55), .b(n123) );
	ao21_6 U106 ( .x(DIFF[8]), .a(A[8]), .b(n87), .c(n88) );
	inv_2 U107 ( .x(n56), .a(n121) );
	nand2i_4 U108 ( .x(n124), .a(A[26]), .b(n57) );
	or3i_5 U109 ( .x(n91), .a(n142), .b(n166), .c(n80) );
	inv_10 U11 ( .x(n79), .a(A[4]) );
	nand2i_4 U110 ( .x(n168), .a(n80), .b(n142) );
	inv_0 U111 ( .x(n162), .a(A[25]) );
	nand3i_1 U112 ( .x(n58), .a(A[7]), .b(n140), .c(n139) );
	inv_10 U113 ( .x(n142), .a(n136) );
	nand2i_4 U115 ( .x(n166), .a(A[9]), .b(n90) );
	inv_5 U116 ( .x(n103), .a(A[15]) );
	nand2i_4 U117 ( .x(n96), .a(n64), .b(n182) );
	nor3_2 U118 ( .x(n115), .a(n54), .b(A[19]), .c(n143) );
	inv_7 U119 ( .x(n178), .a(n54) );
	nor2i_2 U12 ( .x(n138), .a(n148), .b(n149) );
	nor2_3 U120 ( .x(n170), .a(n54), .b(n147) );
	nand2i_1 U121 ( .x(n179), .a(A[15]), .b(n73) );
	nand2_5 U123 ( .x(n61), .a(n106), .b(n103) );
	nand2_6 U124 ( .x(DIFF[23]), .a(n119), .b(n120) );
	nand2_1 U125 ( .x(n70), .a(n146), .b(n142) );
	nand2_6 U126 ( .x(n118), .a(n170), .b(n116) );
	nand2i_4 U127 ( .x(n107), .a(n54), .b(n116) );
	nor2i_3 U128 ( .x(n65), .a(n66), .b(n151) );
	inv_5 U129 ( .x(n153), .a(n65) );
	nor2i_3 U13 ( .x(n137), .a(n138), .b(n70) );
	inv_0 U131 ( .x(n67), .a(A[6]) );
	mux2i_3 U132 ( .x(DIFF[9]), .d0(n141), .sl(A[9]), .d1(n88) );
	nand2_8 U133 ( .x(n111), .a(n146), .b(n142) );
	nor2_1 U134 ( .x(n84), .a(A[2]), .b(A[4]) );
	nor2_1 U135 ( .x(n169), .a(A[2]), .b(A[4]) );
	nand2_0 U136 ( .x(n71), .a(n146), .b(n142) );
	oai22_2 U137 ( .x(DIFF[18]), .a(n112), .b(n71), .c(n113), .d(n114) );
	nand2i_4 U138 ( .x(n143), .a(A[17]), .b(n114) );
	nand3i_3 U139 ( .x(n172), .a(n143), .b(n178), .c(n116) );
	nor2_0 U14 ( .x(n176), .a(A[2]), .b(A[4]) );
	nand2_8 U140 ( .x(n112), .a(n178), .b(n148) );
	inv_0 U141 ( .x(n82), .a(A[5]) );
	oai21_4 U142 ( .x(DIFF[14]), .a(n99), .b(n100), .c(n101) );
	aoai211_4 U143 ( .x(DIFF[20]), .a(n115), .b(n116), .c(n117), .d(n118) );
	nor2i_5 U144 ( .x(n133), .a(n134), .b(n128) );
	nand2_5 U145 ( .x(n128), .a(n156), .b(n157) );
	nor2_5 U146 ( .x(n150), .a(n149), .b(n147) );
	nand2i_4 U147 ( .x(n181), .a(A[2]), .b(n158) );
	nand2i_4 U148 ( .x(n97), .a(A[13]), .b(n116) );
	inv_5 U149 ( .x(n156), .a(n76) );
	nand3i_3 U15 ( .x(n147), .a(A[19]), .b(n117), .c(n148) );
	nand2i_4 U150 ( .x(n129), .a(n157), .b(n76) );
	nand2i_4 U151 ( .x(n77), .a(n159), .b(n126) );
	nand2i_4 U152 ( .x(n122), .a(n163), .b(n119) );
	nand2i_4 U153 ( .x(n120), .a(n164), .b(n153) );
	nand2i_4 U154 ( .x(n98), .a(n165), .b(n96) );
	nand2_6 U155 ( .x(DIFF[26]), .a(n124), .b(n125) );
	nand2_6 U156 ( .x(DIFF[28]), .a(n76), .b(n77) );
	nand2_6 U157 ( .x(DIFF[29]), .a(n128), .b(n129) );
	aoai211_5 U158 ( .x(DIFF[7]), .a(n84), .b(n85), .c(n86), .d(n87) );
	inv_6 U159 ( .x(n94), .a(n93) );
	nor2i_2 U16 ( .x(n177), .a(n109), .b(n54) );
	inv_10 U160 ( .x(n95), .a(A[12]) );
	nand2_8 U161 ( .x(n132), .a(n150), .b(n116) );
	nand2i_6 U162 ( .x(n126), .a(A[27]), .b(n154) );
	nand2i_6 U163 ( .x(n76), .a(A[28]), .b(n155) );
	inv_6 U164 ( .x(n78), .a(n181) );
	inv_6 U165 ( .x(n148), .a(n143) );
	nor2_6 U166 ( .x(n140), .a(A[6]), .b(A[5]) );
	inv_5 U167 ( .x(n81), .a(n80) );
	mux2i_5 U168 ( .x(DIFF[19]), .d0(n137), .sl(n50), .d1(n172) );
	nand2_4 U169 ( .x(n72), .a(n79), .b(n174) );
	mux2_6 U170 ( .x(DIFF[6]), .d0(n60), .sl(n183), .d1(n83) );
	inv_0 U171 ( .x(n183), .a(n67) );
	nand2_1 U172 ( .x(n83), .a(n169), .b(n175) );
	and2_1 U173 ( .x(n60), .a(n176), .b(n175) );
	inv_6 U174 ( .x(n117), .a(A[20]) );
	inv_7 U175 ( .x(n114), .a(A[18]) );
	inv_5 U176 ( .x(n109), .a(A[17]) );
	inv_3 U177 ( .x(n139), .a(A[8]) );
	inv_1 U178 ( .x(n66), .a(A[22]) );
	inv_0 U18 ( .x(n131), .a(A[21]) );
	inv_5 U19 ( .x(n171), .a(n118) );
	inv_5 U20 ( .x(n108), .a(n107) );
	nor2_4 U22 ( .x(n174), .a(A[3]), .b(A[2]) );
	inv_0 U23 ( .x(n161), .a(A[26]) );
	inv_5 U24 ( .x(n154), .a(n124) );
	inv_4 U25 ( .x(n102), .a(n101) );
	oai21_2 U26 ( .x(DIFF[15]), .a(n102), .b(n103), .c(n104) );
	inv_2 U28 ( .x(n99), .a(n97) );
	inv_5 U29 ( .x(n88), .a(n168) );
	ao21_1 U30 ( .x(DIFF[3]), .a(A[3]), .b(A[2]), .c(n78) );
	inv_0 U31 ( .x(DIFF[2]), .a(A[2]) );
	nand2i_2 U32 ( .x(n55), .a(A[25]), .b(n56) );
	inv_4 U33 ( .x(n119), .a(n68) );
	inv_4 U34 ( .x(n113), .a(n110) );
	nor2i_3 U35 ( .x(n68), .a(n164), .b(n153) );
	inv_0 U36 ( .x(n135), .a(A[9]) );
	inv_7 U37 ( .x(n155), .a(n126) );
	oai21_1 U39 ( .x(DIFF[4]), .a(n78), .b(n79), .c(n72) );
	oai21_5 U4 ( .x(DIFF[11]), .a(n92), .b(n75), .c(n93) );
	nand2_3 U40 ( .x(DIFF[13]), .a(n97), .b(n98) );
	inv_7 U41 ( .x(n86), .a(A[7]) );
	exnor2_1 U42 ( .x(DIFF[31]), .a(n133), .b(n167) );
	inv_5 U43 ( .x(n106), .a(A[16]) );
	inv_2 U44 ( .x(n90), .a(A[10]) );
	inv_0 U45 ( .x(n163), .a(A[24]) );
	inv_8 U46 ( .x(n100), .a(A[14]) );
	inv_7 U48 ( .x(n165), .a(A[13]) );
	inv_2 U49 ( .x(n160), .a(A[27]) );
	nand2i_5 U5 ( .x(n151), .a(A[21]), .b(n152) );
	inv_2 U50 ( .x(n159), .a(A[28]) );
	inv_2 U51 ( .x(n157), .a(A[29]) );
	inv_2 U52 ( .x(n167), .a(A[31]) );
	inv_3 U53 ( .x(n75), .a(A[11]) );
	exnor2_5 U54 ( .x(DIFF[30]), .a(n128), .b(n53) );
	buf_1 U55 ( .x(n51), .a(n90) );
	mux2i_3 U56 ( .x(DIFF[21]), .d0(n132), .sl(A[21]), .d1(n171) );
	oai21_5 U57 ( .x(DIFF[16]), .a(n105), .b(n106), .c(n107) );
	nor2_8 U58 ( .x(n145), .a(A[9]), .b(A[10]) );
	nor2_1 U59 ( .x(n175), .a(A[5]), .b(A[3]) );
	inv_10 U6 ( .x(n152), .a(n132) );
	oai21_2 U60 ( .x(DIFF[5]), .a(n81), .b(n82), .c(n83) );
	nand2i_4 U62 ( .x(n141), .a(n72), .b(n142) );
	mux2i_3 U63 ( .x(DIFF[22]), .d0(n130), .sl(n66), .d1(n151) );
	inv_6 U64 ( .x(n105), .a(n104) );
	inv_5 U65 ( .x(n158), .a(A[3]) );
	inv_1 U67 ( .x(n64), .a(n69) );
	inv_1 U68 ( .x(n69), .a(n144) );
	nor3_1 U69 ( .x(n85), .a(A[3]), .b(A[6]), .c(A[5]) );
	nand4i_1 U70 ( .x(n87), .a(A[5]), .b(n173), .c(n174), .d(n79) );
	nor3_5 U71 ( .x(n146), .a(n144), .b(n63), .c(n62) );
	nand2i_3 U72 ( .x(n62), .a(A[2]), .b(n158) );
	nand2_6 U73 ( .x(n101), .a(n73), .b(n116) );
	nand2_6 U74 ( .x(n59), .a(n165), .b(n100) );
	inv_7 U75 ( .x(n73), .a(n59) );
	and4i_1 U76 ( .x(n52), .a(n151), .b(n163), .c(n164), .d(n66) );
	inv_3 U77 ( .x(n121), .a(n52) );
	inv_2 U78 ( .x(n164), .a(A[23]) );
	nor2_3 U79 ( .x(n180), .a(n72), .b(n166) );
	inv_2 U8 ( .x(n50), .a(A[19]) );
	oai21_5 U80 ( .x(DIFF[12]), .a(n94), .b(n95), .c(n96) );
	inv_6 U81 ( .x(n63), .a(n79) );
	nand2_3 U82 ( .x(n80), .a(n79), .b(n174) );
	nand2_6 U83 ( .x(DIFF[27]), .a(n126), .b(n127) );
	nand3_3 U84 ( .x(n93), .a(n142), .b(n75), .c(n180) );
	nand3i_5 U85 ( .x(n144), .a(A[11]), .b(n95), .c(n145) );
	nand3_4 U86 ( .x(n136), .a(n86), .b(n139), .c(n140) );
	nand2i_3 U88 ( .x(n104), .a(n179), .b(n116) );
	inv_2 U89 ( .x(n53), .a(n134) );
	nand2_6 U9 ( .x(DIFF[24]), .a(n121), .b(n122) );
	inv_2 U90 ( .x(n134), .a(A[30]) );
	nor2_2 U91 ( .x(n173), .a(A[7]), .b(A[6]) );
	inv_6 U92 ( .x(n92), .a(n91) );
	nand2i_6 U93 ( .x(n149), .a(n61), .b(n73) );
	nand2i_6 U94 ( .x(n54), .a(n61), .b(n73) );
	inv_16 U95 ( .x(n116), .a(n111) );
	inv_4 U96 ( .x(n182), .a(n141) );
	oai21_2 U97 ( .x(DIFF[10]), .a(n89), .b(n51), .c(n91) );
	nor3i_2 U98 ( .x(n89), .a(n135), .b(n72), .c(n58) );
	oai21_4 U99 ( .x(DIFF[17]), .a(n108), .b(n109), .c(n110) );

endmodule


module ID_DW01_sub_32_1_test_1 (  A, B, CI, DIFF, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] DIFF;

wire A_0, A_1, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
	n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
	n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
	n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
	n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
	n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
	n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n51, n52,
	n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
	n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
	n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
	n95, n96, n97, n98, n99;

	assign A_1 = A[1];
	assign A_0 = A[0];
	assign DIFF[1] = A_1;
	assign DIFF[0] = A_0;

	nor2_0 U10 ( .x(n166), .a(A[2]), .b(A[3]) );
	nor2_2 U100 ( .x(n167), .a(A[2]), .b(A[3]) );
	and4i_4 U101 ( .x(n58), .a(n59), .b(n154), .c(n155), .d(n156) );
	inv_4 U102 ( .x(n78), .a(n58) );
	inv_2 U103 ( .x(n59), .a(n157) );
	ao21_4 U104 ( .x(DIFF[14]), .a(n83), .b(A[14]), .c(n60) );
	nor2_1 U105 ( .x(n161), .a(A[2]), .b(A[3]) );
	nor2_5 U106 ( .x(n60), .a(n129), .b(n79) );
	inv_10 U107 ( .x(n134), .a(n79) );
	nor2_1 U108 ( .x(n131), .a(A[6]), .b(A[10]) );
	aoi21_1 U109 ( .x(n62), .a(n132), .b(n166), .c(n128) );
	inv_0 U11 ( .x(n136), .a(n54) );
	nand2i_0 U110 ( .x(n174), .a(A[15]), .b(n173) );
	nand3i_1 U111 ( .x(n135), .a(A[15]), .b(n94), .c(n168) );
	inv_0 U112 ( .x(n151), .a(A[15]) );
	nor2_0 U113 ( .x(n175), .a(A[15]), .b(A[16]) );
	nand2_1 U114 ( .x(n92), .a(A[17]), .b(n90) );
	inv_2 U116 ( .x(DIFF[2]), .a(A[2]) );
	nand2_6 U117 ( .x(DIFF[27]), .a(n116), .b(n117) );
	nand2i_6 U118 ( .x(n116), .a(A[27]), .b(n143) );
	nor2_0 U119 ( .x(n170), .a(A[21]), .b(A[20]) );
	nand2i_0 U12 ( .x(n140), .a(A[25]), .b(n114) );
	ao21_1 U120 ( .x(DIFF[3]), .a(A[3]), .b(A[2]), .c(n68) );
	and4i_3 U121 ( .x(n65), .a(n66), .b(n131), .c(n132), .d(n133) );
	nor2_0 U122 ( .x(n125), .a(A[5]), .b(A[6]) );
	nand3i_1 U123 ( .x(n129), .a(A[13]), .b(n85), .c(n130) );
	inv_0 U124 ( .x(n153), .a(A[13]) );
	nand2i_2 U125 ( .x(n70), .a(n63), .b(n161) );
	mux2i_2 U126 ( .x(DIFF[11]), .d0(n162), .sl(A[11]), .d1(n134) );
	nor2_0 U128 ( .x(n173), .a(A[17]), .b(A[16]) );
	inv_0 U129 ( .x(n158), .a(A[10]) );
	oai21_2 U13 ( .x(DIFF[18]), .a(n93), .b(n94), .c(n64) );
	nand2_1 U130 ( .x(n67), .a(n127), .b(n69) );
	inv_2 U131 ( .x(n155), .a(n67) );
	inv_0 U132 ( .x(n176), .a(A[11]) );
	nand2i_2 U133 ( .x(n162), .a(A[10]), .b(n58) );
	nand4i_1 U134 ( .x(n72), .a(A[7]), .b(n164), .c(n165), .d(n69) );
	oai21_1 U135 ( .x(n82), .a(A[11]), .b(n79), .c(A[12]) );
	nand2i_0 U136 ( .x(n152), .a(A[12]), .b(n176) );
	nor2_0 U137 ( .x(n165), .a(A[6]), .b(A[5]) );
	oai21_4 U138 ( .x(DIFF[4]), .a(n68), .b(n69), .c(n70) );
	oai21_4 U139 ( .x(DIFF[9]), .a(n76), .b(n77), .c(n78) );
	inv_2 U14 ( .x(n93), .a(n91) );
	oai21_4 U140 ( .x(DIFF[20]), .a(n98), .b(n99), .c(n100) );
	oai21_4 U141 ( .x(DIFF[21]), .a(n101), .b(n102), .c(n103) );
	oai21_4 U142 ( .x(DIFF[22]), .a(n104), .b(n105), .c(n106) );
	oai21_4 U143 ( .x(DIFF[24]), .a(n109), .b(n110), .c(n111) );
	nand2i_4 U144 ( .x(n74), .a(n163), .b(n178) );
	nand2i_4 U145 ( .x(n75), .a(n51), .b(n72) );
	nand2i_4 U146 ( .x(n86), .a(A[15]), .b(n60) );
	inv_5 U147 ( .x(n88), .a(n86) );
	nand2i_4 U148 ( .x(n91), .a(n174), .b(n60) );
	nand2i_4 U149 ( .x(n100), .a(n172), .b(n137) );
	nand2_2 U15 ( .x(DIFF[17]), .a(n91), .b(n92) );
	nand2i_4 U150 ( .x(n103), .a(n171), .b(n137) );
	nand2i_4 U151 ( .x(n107), .a(A[23]), .b(n139) );
	nand2i_4 U152 ( .x(n113), .a(n148), .b(n111) );
	nand2i_4 U153 ( .x(n108), .a(n149), .b(n106) );
	nand2i_4 U154 ( .x(n84), .a(n153), .b(n81) );
	nand2i_4 U155 ( .x(n80), .a(n158), .b(n78) );
	nand2_5 U156 ( .x(DIFF[23]), .a(n107), .b(n108) );
	nand2_5 U157 ( .x(DIFF[25]), .a(n112), .b(n113) );
	oai21_5 U158 ( .x(DIFF[28]), .a(n118), .b(n119), .c(n120) );
	exnor2_5 U159 ( .x(DIFF[30]), .a(n160), .b(n124) );
	nand2i_2 U16 ( .x(n138), .a(A[23]), .b(n110) );
	nand2i_6 U160 ( .x(n81), .a(n152), .b(n134) );
	nand2i_6 U161 ( .x(n111), .a(n138), .b(n139) );
	nand2i_6 U162 ( .x(n120), .a(n142), .b(n143) );
	mux2i_1 U163 ( .x(n55), .d0(n56), .sl(A[5]), .d1(n70) );
	inv_0 U164 ( .x(n99), .a(A[20]) );
	inv_0 U165 ( .x(n94), .a(A[18]) );
	inv_2 U166 ( .x(n110), .a(A[24]) );
	nor2_1 U167 ( .x(n168), .a(A[17]), .b(A[16]) );
	inv_4 U168 ( .x(n51), .a(A[8]) );
	nand2i_1 U169 ( .x(n163), .a(A[8]), .b(n127) );
	nand2i_2 U17 ( .x(n87), .a(n151), .b(n61) );
	inv_5 U170 ( .x(n105), .a(A[22]) );
	nand2_3 U18 ( .x(DIFF[8]), .a(n74), .b(n75) );
	inv_4 U19 ( .x(n76), .a(n74) );
	nand2i_0 U20 ( .x(n171), .a(A[19]), .b(n170) );
	nand2i_0 U21 ( .x(n172), .a(A[19]), .b(n99) );
	nand2i_2 U23 ( .x(n122), .a(n146), .b(n120) );
	nand2i_2 U24 ( .x(n177), .a(A[2]), .b(n145) );
	inv_5 U25 ( .x(n179), .a(n81) );
	nand2i_2 U26 ( .x(n117), .a(n147), .b(n115) );
	inv_2 U27 ( .x(n118), .a(n116) );
	nand2_2 U28 ( .x(DIFF[7]), .a(n72), .b(n73) );
	nand2i_2 U29 ( .x(n96), .a(A[19]), .b(n137) );
	nand2_2 U30 ( .x(DIFF[19]), .a(n96), .b(n97) );
	nand2i_2 U31 ( .x(n97), .a(n150), .b(n64) );
	inv_2 U32 ( .x(n98), .a(n96) );
	inv_5 U33 ( .x(n141), .a(n111) );
	inv_7 U34 ( .x(n139), .a(n106) );
	nand2_2 U35 ( .x(DIFF[15]), .a(n86), .b(n87) );
	inv_4 U36 ( .x(n68), .a(n177) );
	inv_2 U37 ( .x(n101), .a(n100) );
	inv_0 U38 ( .x(n85), .a(A[14]) );
	inv_2 U39 ( .x(n109), .a(n107) );
	nand2_2 U4 ( .x(DIFF[10]), .a(n80), .b(n79) );
	inv_2 U40 ( .x(n104), .a(n103) );
	nand2_2 U41 ( .x(DIFF[29]), .a(n121), .b(n122) );
	inv_3 U42 ( .x(n127), .a(A[7]) );
	exnor2_1 U43 ( .x(DIFF[31]), .a(n123), .b(n159) );
	nor2i_1 U44 ( .x(n123), .a(n124), .b(n121) );
	inv_2 U45 ( .x(n144), .a(n120) );
	nand2i_2 U46 ( .x(n121), .a(A[29]), .b(n144) );
	inv_2 U47 ( .x(n160), .a(n121) );
	inv_0 U48 ( .x(n114), .a(A[26]) );
	inv_0 U5 ( .x(n150), .a(A[19]) );
	inv_0 U51 ( .x(n148), .a(A[25]) );
	inv_0 U52 ( .x(n102), .a(A[21]) );
	inv_2 U54 ( .x(n149), .a(A[23]) );
	inv_2 U55 ( .x(n147), .a(A[27]) );
	inv_2 U56 ( .x(n119), .a(A[28]) );
	inv_2 U57 ( .x(n146), .a(A[29]) );
	inv_2 U58 ( .x(n124), .a(A[30]) );
	inv_2 U59 ( .x(n159), .a(A[31]) );
	nand2i_2 U6 ( .x(n142), .a(A[27]), .b(n119) );
	inv_4 U60 ( .x(n63), .a(n69) );
	ao21_4 U61 ( .x(DIFF[26]), .a(n112), .b(A[26]), .c(n143) );
	inv_2 U62 ( .x(n61), .a(n60) );
	nand2i_2 U63 ( .x(n64), .a(n135), .b(n60) );
	nand2i_3 U64 ( .x(n95), .a(n135), .b(n60) );
	nand3i_2 U65 ( .x(n90), .a(n129), .b(n175), .c(n134) );
	inv_8 U66 ( .x(n79), .a(n65) );
	oai21_5 U67 ( .x(DIFF[16]), .a(n88), .b(n89), .c(n90) );
	nor2_2 U68 ( .x(n132), .a(A[4]), .b(A[5]) );
	inv_5 U7 ( .x(n69), .a(A[4]) );
	nor2_0 U70 ( .x(n154), .a(A[5]), .b(A[6]) );
	inv_5 U71 ( .x(n143), .a(n115) );
	nand2i_5 U72 ( .x(n112), .a(A[25]), .b(n141) );
	nand2_8 U73 ( .x(DIFF[13]), .a(n83), .b(n84) );
	nand2i_5 U74 ( .x(n83), .a(A[13]), .b(n179) );
	and2_2 U75 ( .x(n156), .a(n77), .b(n51) );
	inv_4 U76 ( .x(n77), .a(A[9]) );
	nor2_5 U77 ( .x(n133), .a(A[2]), .b(A[3]) );
	inv_2 U78 ( .x(n57), .a(n63) );
	inv_3 U79 ( .x(n145), .a(A[3]) );
	nand3_1 U8 ( .x(n71), .a(n69), .b(n125), .c(n126) );
	nor2_1 U80 ( .x(n157), .a(A[2]), .b(A[3]) );
	nor2_1 U81 ( .x(n164), .a(A[2]), .b(A[3]) );
	nand2i_2 U82 ( .x(n73), .a(n127), .b(n71) );
	inv_4 U83 ( .x(n178), .a(n71) );
	inv_0 U84 ( .x(n89), .a(A[16]) );
	or2_6 U85 ( .x(DIFF[6]), .a(n178), .b(n62) );
	nand3_1 U86 ( .x(n66), .a(n127), .b(n51), .c(n77) );
	nand2_3 U87 ( .x(DIFF[12]), .a(n81), .b(n82) );
	nand4i_1 U88 ( .x(n115), .a(n140), .b(n52), .c(n137), .d(n54) );
	inv_2 U89 ( .x(n52), .a(n138) );
	inv_0 U9 ( .x(n128), .a(A[6]) );
	inv_7 U90 ( .x(n137), .a(n95) );
	nor2_3 U91 ( .x(n126), .a(A[2]), .b(A[3]) );
	nand2_8 U92 ( .x(n106), .a(n53), .b(n137) );
	inv_2 U93 ( .x(n53), .a(n136) );
	and3_1 U94 ( .x(n54), .a(n150), .b(n105), .c(n169) );
	nor2_0 U95 ( .x(n169), .a(A[21]), .b(A[20]) );
	nor2_1 U97 ( .x(n130), .a(A[12]), .b(A[11]) );
	inv_5 U98 ( .x(DIFF[5]), .a(n55) );
	and2_5 U99 ( .x(n56), .a(n57), .b(n167) );

endmodule


module ID_DW01_add_32_0_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
	n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
	n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
	n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
	n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
	n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
	n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
	n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
	n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
	n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
	n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
	n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
	n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399,
	n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
	n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423,
	n424, n425, n426, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
	n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
	n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
	n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99;


	nand2_2 U10 ( .x(n353), .a(B[30]), .b(n70) );
	inv_2 U100 ( .x(n320), .a(n99) );
	nand2i_2 U101 ( .x(n325), .a(n320), .b(n321) );
	nand2i_2 U102 ( .x(n330), .a(n173), .b(n413) );
	nand2_0 U103 ( .x(n172), .a(A[10]), .b(B[10]) );
	inv_2 U104 ( .x(n291), .a(n137) );
	nand2i_2 U105 ( .x(n369), .a(n370), .b(n371) );
	nand2i_3 U106 ( .x(n249), .a(A[15]), .b(n237) );
	nand2_0 U107 ( .x(n158), .a(B[15]), .b(A[15]) );
	nand2i_2 U108 ( .x(n397), .a(A[14]), .b(n238) );
	nor2i_1 U109 ( .x(n180), .a(n181), .b(n182) );
	nand2i_2 U11 ( .x(n279), .a(n70), .b(n408) );
	inv_5 U110 ( .x(n182), .a(n414) );
	nand2i_2 U111 ( .x(n327), .a(B[10]), .b(n243) );
	inv_2 U112 ( .x(n329), .a(n172) );
	nand2_2 U113 ( .x(n96), .a(A[8]), .b(B[8]) );
	ao21_1 U114 ( .x(n398), .a(n233), .b(n232), .c(n96) );
	nand2i_2 U115 ( .x(n245), .a(B[8]), .b(n231) );
	nand2i_2 U116 ( .x(n244), .a(n190), .b(n245) );
	nand2i_2 U117 ( .x(n384), .a(B[3]), .b(n227) );
	inv_1 U118 ( .x(n227), .a(A[3]) );
	nand2_0 U119 ( .x(n121), .a(A[3]), .b(B[3]) );
	nand2_2 U12 ( .x(n408), .a(B[27]), .b(B[26]) );
	inv_2 U120 ( .x(n226), .a(B[2]) );
	inv_5 U121 ( .x(n396), .a(n395) );
	nand2_2 U122 ( .x(n393), .a(B[25]), .b(n70) );
	inv_5 U123 ( .x(n270), .a(B[25]) );
	inv_2 U124 ( .x(n272), .a(B[24]) );
	nand2i_2 U125 ( .x(n394), .a(B[24]), .b(n273) );
	nand2_2 U126 ( .x(n371), .a(n286), .b(n287) );
	inv_2 U127 ( .x(n367), .a(n371) );
	inv_2 U128 ( .x(n368), .a(n134) );
	nor2i_1 U129 ( .x(n366), .a(n139), .b(n368) );
	nand2_0 U13 ( .x(n347), .a(B[27]), .b(B[26]) );
	nor2i_1 U130 ( .x(n83), .a(n366), .b(n367) );
	nand2_2 U131 ( .x(n364), .a(n365), .b(n263) );
	nand2i_2 U132 ( .x(n262), .a(A[21]), .b(n274) );
	inv_2 U133 ( .x(n274), .a(B[21]) );
	nand2_2 U134 ( .x(n137), .a(B[21]), .b(A[21]) );
	oai31_2 U135 ( .x(n346), .a(n339), .b(n182), .c(n338), .d(n344) );
	inv_7 U136 ( .x(n334), .a(n248) );
	inv_5 U137 ( .x(n335), .a(n246) );
	nand2_2 U138 ( .x(n333), .a(n334), .b(n335) );
	inv_2 U139 ( .x(n235), .a(A[20]) );
	nor2_1 U14 ( .x(n200), .a(A[22]), .b(B[22]) );
	aoi21_1 U140 ( .x(n341), .a(n323), .b(n342), .c(n343) );
	inv_2 U141 ( .x(n343), .a(n146) );
	inv_5 U142 ( .x(n332), .a(n239) );
	inv_2 U143 ( .x(n254), .a(B[17]) );
	inv_2 U144 ( .x(n380), .a(n152) );
	nand2_2 U145 ( .x(n152), .a(n62), .b(A[17]) );
	inv_1 U146 ( .x(n316), .a(n412) );
	inv_2 U147 ( .x(n258), .a(A[18]) );
	nor2i_1 U148 ( .x(n315), .a(n152), .b(n258) );
	nor2i_1 U149 ( .x(n314), .a(n315), .b(n316) );
	nor2_4 U15 ( .x(n265), .a(n199), .b(n200) );
	inv_2 U150 ( .x(n271), .a(B[23]) );
	inv_2 U151 ( .x(n370), .a(n139) );
	nand2_2 U152 ( .x(n139), .a(A[23]), .b(B[23]) );
	inv_2 U153 ( .x(n365), .a(n289) );
	nand2i_2 U154 ( .x(n289), .a(n136), .b(n262) );
	inv_2 U155 ( .x(n136), .a(n293) );
	nor2_1 U156 ( .x(n135), .a(n136), .b(n137) );
	nor2i_1 U157 ( .x(n372), .a(n373), .b(n135) );
	inv_2 U158 ( .x(n234), .a(B[30]) );
	nand2i_0 U159 ( .x(n355), .a(n125), .b(n351) );
	nand2i_4 U16 ( .x(n264), .a(B[24]), .b(n273) );
	inv_5 U160 ( .x(n351), .a(n277) );
	nor2i_1 U161 ( .x(n356), .a(n357), .b(n358) );
	inv_2 U162 ( .x(n357), .a(n282) );
	inv_2 U163 ( .x(n358), .a(n124) );
	inv_2 U164 ( .x(n406), .a(n285) );
	oai211_1 U165 ( .x(n119), .a(n348), .b(n196), .c(n281), .d(n354) );
	nand2_2 U166 ( .x(n108), .a(B[4]), .b(A[4]) );
	inv_2 U167 ( .x(n225), .a(B[4]) );
	inv_2 U168 ( .x(n165), .a(n181) );
	nand2_2 U169 ( .x(n164), .a(A[13]), .b(B[13]) );
	nand2_0 U17 ( .x(n283), .a(B[28]), .b(n70) );
	nand2i_0 U170 ( .x(n116), .a(n378), .b(n167) );
	nor2_0 U171 ( .x(n115), .a(n247), .b(n170) );
	inv_4 U172 ( .x(n247), .a(n420) );
	nand2i_2 U173 ( .x(n111), .a(B[11]), .b(n252) );
	exor2_1 U174 ( .x(n213), .a(B[27]), .b(n70) );
	inv_2 U175 ( .x(n129), .a(n131) );
	exor2_1 U176 ( .x(SUM[7]), .a(n205), .b(n98) );
	ao21_1 U177 ( .x(n205), .a(n322), .b(n391), .c(n390) );
	inv_2 U178 ( .x(n390), .a(n102) );
	nor2i_1 U179 ( .x(n98), .a(n99), .b(n100) );
	inv_5 U18 ( .x(n269), .a(B[28]) );
	inv_2 U180 ( .x(n100), .a(n382) );
	aoi21_1 U181 ( .x(n85), .a(n86), .b(n69), .c(n88) );
	exnor2_1 U182 ( .x(n308), .a(B[29]), .b(n70) );
	inv_2 U183 ( .x(n125), .a(n381) );
	nor2i_1 U184 ( .x(n123), .a(n124), .b(n125) );
	nor2i_1 U185 ( .x(n130), .a(n131), .b(n132) );
	inv_2 U186 ( .x(n132), .a(n127) );
	exnor2_1 U187 ( .x(SUM[8]), .a(n51), .b(n95) );
	nor2i_1 U188 ( .x(n95), .a(n96), .b(n97) );
	exnor2_1 U189 ( .x(SUM[12]), .a(n110), .b(n166) );
	nor2i_1 U19 ( .x(n192), .a(n137), .b(n193) );
	inv_2 U190 ( .x(n113), .a(n169) );
	nor2i_1 U191 ( .x(n166), .a(n167), .b(n109) );
	exor2_1 U192 ( .x(SUM[16]), .a(n219), .b(n154) );
	nand2i_2 U193 ( .x(n219), .a(n295), .b(n401) );
	nor2i_1 U194 ( .x(n154), .a(n155), .b(n156) );
	nand2i_2 U195 ( .x(n78), .a(n52), .b(n203) );
	inv_2 U196 ( .x(n422), .a(n421) );
	mux2i_1 U197 ( .x(n77), .d0(n422), .sl(A[19]), .d1(n305) );
	nand2_2 U198 ( .x(SUM[19]), .a(n77), .b(n78) );
	exor2_1 U199 ( .x(SUM[20]), .a(n216), .b(n145) );
	nand2i_2 U20 ( .x(n301), .a(A[18]), .b(n259) );
	nand2i_2 U200 ( .x(n216), .a(n376), .b(n410) );
	nor2i_1 U201 ( .x(n145), .a(n146), .b(n147) );
	inv_5 U202 ( .x(n147), .a(n342) );
	exor2_1 U203 ( .x(SUM[9]), .a(n204), .b(n93) );
	oai21_1 U204 ( .x(n204), .a(n51), .b(n97), .c(n96) );
	inv_2 U205 ( .x(n97), .a(n245) );
	nor2i_1 U206 ( .x(n93), .a(n94), .b(n92) );
	inv_2 U207 ( .x(n156), .a(n241) );
	exor2_1 U208 ( .x(SUM[17]), .a(n66), .b(n151) );
	nor2i_1 U209 ( .x(SUM[0]), .a(n73), .b(n74) );
	nor3_0 U21 ( .x(n299), .a(n153), .b(n156), .c(n240) );
	nand2_2 U210 ( .x(n73), .a(B[0]), .b(A[0]) );
	nor2i_1 U211 ( .x(n168), .a(n169), .b(n170) );
	inv_2 U212 ( .x(n170), .a(n111) );
	exor2_1 U213 ( .x(SUM[24]), .a(n214), .b(n133) );
	nand2i_2 U214 ( .x(n214), .a(n369), .b(n82) );
	nor2i_1 U215 ( .x(n133), .a(n134), .b(n84) );
	inv_2 U216 ( .x(n159), .a(n249) );
	exor2_1 U217 ( .x(SUM[15]), .a(n220), .b(n157) );
	inv_2 U218 ( .x(n400), .a(n221) );
	nand2i_2 U219 ( .x(n221), .a(n180), .b(n399) );
	ao221_2 U22 ( .x(n256), .a(n254), .b(n253), .c(n155), .d(n257), .e(n240) );
	ao21_3 U220 ( .x(n208), .a(n384), .b(n212), .c(n59) );
	nor2i_1 U221 ( .x(n107), .a(n108), .b(n91) );
	exor2_1 U222 ( .x(SUM[10]), .a(n222), .b(n171) );
	oai211_1 U223 ( .x(n222), .a(n51), .b(n244), .c(n398), .d(n94) );
	nor2i_1 U224 ( .x(n171), .a(n172), .b(n173) );
	inv_2 U225 ( .x(n173), .a(n327) );
	exor2_1 U226 ( .x(SUM[3]), .a(n212), .b(n120) );
	inv_2 U227 ( .x(n387), .a(n149) );
	nor2i_1 U228 ( .x(n120), .a(n121), .b(n122) );
	inv_2 U229 ( .x(n122), .a(n384) );
	nand2i_0 U23 ( .x(n297), .a(n298), .b(n256) );
	exor2_1 U230 ( .x(SUM[2]), .a(n426), .b(n148) );
	oai21_2 U231 ( .x(n217), .a(n176), .b(n73), .c(n175) );
	nor2i_1 U232 ( .x(n148), .a(n149), .b(n150) );
	inv_2 U233 ( .x(n150), .a(n385) );
	nand2i_2 U234 ( .x(n303), .a(n396), .b(n393) );
	inv_2 U235 ( .x(n84), .a(n394) );
	aoi21_1 U236 ( .x(n81), .a(n82), .b(n83), .c(n84) );
	exnor2_1 U237 ( .x(SUM[25]), .a(n81), .b(n303) );
	inv_2 U238 ( .x(n142), .a(n262) );
	nor2i_1 U239 ( .x(n141), .a(n137), .b(n142) );
	ao21_2 U24 ( .x(n229), .a(n224), .b(n223), .c(n106) );
	exor2_1 U240 ( .x(SUM[21]), .a(n69), .b(n141) );
	ao21_1 U241 ( .x(n76), .a(n152), .b(n412), .c(n301) );
	exor2_1 U242 ( .x(SUM[23]), .a(n215), .b(n138) );
	nor2i_1 U243 ( .x(n138), .a(n139), .b(n140) );
	exnor2_1 U244 ( .x(SUM[1]), .a(n174), .b(n73) );
	nor2i_0 U245 ( .x(n174), .a(n175), .b(n176) );
	inv_5 U247 ( .x(n106), .a(n389) );
	nor2i_0 U248 ( .x(n104), .a(n105), .b(n106) );
	inv_2 U249 ( .x(n383), .a(n108) );
	nand2_1 U25 ( .x(n94), .a(A[9]), .b(B[9]) );
	inv_0 U250 ( .x(n250), .a(A[12]) );
	aoi21_1 U251 ( .x(n51), .a(n317), .b(n392), .c(n319) );
	exnor2_3 U253 ( .x(n304), .a(n290), .b(n53) );
	inv_2 U254 ( .x(n53), .a(n195) );
	inv_2 U255 ( .x(n195), .a(B[22]) );
	inv_2 U256 ( .x(n71), .a(A[31]) );
	inv_2 U257 ( .x(n72), .a(A[31]) );
	buf_1 U258 ( .x(n54), .a(n63) );
	nand2_1 U259 ( .x(n146), .a(B[20]), .b(A[20]) );
	nor2_1 U26 ( .x(n191), .a(B[9]), .b(A[9]) );
	inv_0 U260 ( .x(n178), .a(B[5]) );
	exnor2_3 U261 ( .x(SUM[27]), .a(n126), .b(n213) );
	aoi21_3 U262 ( .x(n126), .a(n127), .b(n128), .c(n129) );
	inv_2 U263 ( .x(n407), .a(n128) );
	exor2_1 U264 ( .x(SUM[26]), .a(n128), .b(n130) );
	inv_0 U265 ( .x(n55), .a(n112) );
	inv_2 U266 ( .x(n56), .a(n55) );
	aoi31_6 U267 ( .x(n186), .a(n63), .b(n108), .c(n187), .d(n188) );
	nand2i_2 U268 ( .x(n293), .a(A[22]), .b(n195) );
	nand2_0 U269 ( .x(n373), .a(A[22]), .b(B[22]) );
	oai21_1 U27 ( .x(n413), .a(n191), .b(n96), .c(n94) );
	nor2i_2 U270 ( .x(n193), .a(A[22]), .b(n195) );
	and3i_1 U271 ( .x(n57), .a(n346), .b(n68), .c(n403) );
	oa31_4 U272 ( .x(n68), .a(n239), .b(n147), .c(n296), .d(n341) );
	nand3i_0 U273 ( .x(n392), .a(n179), .b(n108), .c(n63) );
	nand3i_0 U274 ( .x(n391), .a(n177), .b(n108), .c(n54) );
	oai21_5 U275 ( .x(n63), .a(A[4]), .b(n64), .c(n208) );
	nand2_1 U276 ( .x(n202), .a(B[18]), .b(A[18]) );
	nor2i_0 U277 ( .x(n160), .a(n161), .b(n162) );
	oai21_1 U278 ( .x(n220), .a(n162), .b(n400), .c(n161) );
	mux2i_2 U279 ( .x(n75), .d0(n306), .sl(n58), .d1(n314) );
	nand2i_2 U28 ( .x(n292), .a(n142), .b(n87) );
	inv_2 U280 ( .x(n58), .a(n61) );
	inv_2 U281 ( .x(n87), .a(n57) );
	nand2i_4 U282 ( .x(n420), .a(B[12]), .b(n250) );
	nor2_0 U283 ( .x(n109), .a(B[12]), .b(A[12]) );
	inv_2 U284 ( .x(n238), .a(B[14]) );
	nand2_2 U285 ( .x(n161), .a(B[14]), .b(A[14]) );
	exnor2_5 U286 ( .x(SUM[31]), .a(n117), .b(n209) );
	aoai211_1 U287 ( .x(n206), .a(n108), .b(n54), .c(n106), .d(n105) );
	inv_2 U288 ( .x(n59), .a(n121) );
	inv_0 U289 ( .x(n60), .a(A[11]) );
	inv_4 U29 ( .x(n345), .a(n256) );
	and3i_3 U290 ( .x(n67), .a(n346), .b(n68), .c(n403) );
	mux2i_1 U291 ( .x(SUM[29]), .d0(n123), .sl(n85), .d1(n308) );
	exor2_1 U292 ( .x(SUM[4]), .a(n424), .b(n107) );
	ao21_1 U293 ( .x(n207), .a(n388), .b(n424), .c(n383) );
	inv_0 U294 ( .x(n61), .a(n259) );
	buf_1 U295 ( .x(n62), .a(B[17]) );
	nand2i_4 U296 ( .x(n412), .a(n153), .b(n218) );
	inv_2 U297 ( .x(n153), .a(n402) );
	oai21_4 U298 ( .x(n379), .a(n186), .b(n325), .c(n326) );
	nand2i_3 U299 ( .x(n382), .a(A[7]), .b(n224) );
	inv_4 U30 ( .x(n259), .a(B[18]) );
	inv_0 U300 ( .x(n223), .a(A[7]) );
	inv_0 U301 ( .x(n231), .a(A[8]) );
	inv_2 U302 ( .x(n64), .a(n225) );
	exor2_1 U303 ( .x(SUM[11]), .a(n56), .b(n168) );
	aoi21_1 U304 ( .x(n110), .a(n111), .b(n56), .c(n113) );
	aoi21_1 U305 ( .x(n114), .a(n115), .b(n56), .c(n116) );
	nand2i_2 U306 ( .x(n399), .a(n246), .b(n112) );
	nand2i_4 U307 ( .x(n112), .a(n374), .b(n379) );
	inv_0 U308 ( .x(n243), .a(A[10]) );
	nand2_2 U31 ( .x(n257), .a(B[17]), .b(A[17]) );
	inv_2 U310 ( .x(n65), .a(n211) );
	exor2_1 U312 ( .x(n211), .a(B[30]), .b(n70) );
	aoai211_1 U313 ( .x(n66), .a(n411), .b(n401), .c(n156), .d(n155) );
	nand2i_2 U314 ( .x(n419), .a(A[24]), .b(n272) );
	nand2_1 U315 ( .x(n276), .a(A[24]), .b(B[24]) );
	nand2_0 U316 ( .x(n134), .a(A[24]), .b(B[24]) );
	inv_0 U317 ( .x(n273), .a(A[24]) );
	nand2_2 U318 ( .x(n187), .a(A[5]), .b(B[5]) );
	nor2i_0 U319 ( .x(n179), .a(A[5]), .b(n178) );
	inv_2 U32 ( .x(n253), .a(A[17]) );
	nor2i_0 U320 ( .x(n177), .a(A[5]), .b(n178) );
	nand2_0 U321 ( .x(n105), .a(A[5]), .b(B[5]) );
	nor2_0 U322 ( .x(n74), .a(A[0]), .b(B[0]) );
	inv_0 U323 ( .x(n251), .a(A[13]) );
	inv_0 U324 ( .x(n233), .a(A[9]) );
	nor2_1 U325 ( .x(n190), .a(B[9]), .b(A[9]) );
	nor2_0 U326 ( .x(n92), .a(B[9]), .b(A[9]) );
	inv_10 U327 ( .x(n69), .a(n67) );
	or3i_5 U328 ( .x(n403), .a(n415), .b(n333), .c(n331) );
	nand3i_2 U329 ( .x(n321), .a(n100), .b(A[6]), .c(B[6]) );
	inv_2 U33 ( .x(n298), .a(n202) );
	nand2_0 U330 ( .x(n102), .a(A[6]), .b(B[6]) );
	inv_0 U331 ( .x(n252), .a(A[11]) );
	nand2i_0 U332 ( .x(n388), .a(A[4]), .b(n225) );
	nor2_0 U333 ( .x(n91), .a(A[4]), .b(B[4]) );
	nand2i_2 U334 ( .x(n385), .a(A[2]), .b(n226) );
	nand2_2 U335 ( .x(n149), .a(B[2]), .b(A[2]) );
	nand2_2 U336 ( .x(n175), .a(A[1]), .b(B[1]) );
	inv_16 U337 ( .x(n70), .a(n71) );
	nor2i_5 U338 ( .x(n101), .a(n102), .b(n103) );
	aoi21_3 U339 ( .x(n117), .a(n118), .b(n69), .c(n119) );
	nor3_2 U34 ( .x(n201), .a(n147), .b(n202), .c(n203) );
	nor2i_5 U340 ( .x(n151), .a(n152), .b(n153) );
	nor2i_5 U341 ( .x(n163), .a(n164), .b(n165) );
	nor2_5 U342 ( .x(n189), .a(A[19]), .b(B[19]) );
	nor2_5 U343 ( .x(n194), .a(A[17]), .b(B[17]) );
	nor2_5 U344 ( .x(n196), .a(n197), .b(n198) );
	exor2_3 U345 ( .x(SUM[6]), .a(n206), .b(n101) );
	exor2_3 U346 ( .x(SUM[5]), .a(n207), .b(n104) );
	exor2_3 U347 ( .x(SUM[14]), .a(n221), .b(n160) );
	exnor2_5 U348 ( .x(SUM[13]), .a(n114), .b(n163) );
	inv_6 U349 ( .x(n237), .a(B[15]) );
	nand2_2 U35 ( .x(n167), .a(A[12]), .b(B[12]) );
	nand3i_5 U350 ( .x(n239), .a(n240), .b(n241), .c(n242) );
	ao21_4 U351 ( .x(n266), .a(n72), .b(n234), .c(n125) );
	oai211_4 U352 ( .x(n198), .a(n71), .b(n270), .c(n139), .d(n276) );
	nand2i_4 U353 ( .x(n277), .a(n278), .b(n279) );
	nand2i_4 U354 ( .x(n290), .a(n291), .b(n292) );
	exnor2_3 U355 ( .x(n306), .a(A[18]), .b(n307) );
	nor2i_5 U356 ( .x(n309), .a(n310), .b(n284) );
	nand2i_4 U358 ( .x(n188), .a(n103), .b(n324) );
	nor2i_5 U359 ( .x(n326), .a(n327), .b(n244) );
	nand2i_2 U36 ( .x(n328), .a(n329), .b(n330) );
	nand2i_4 U360 ( .x(n331), .a(n147), .b(n332) );
	nor2i_5 U361 ( .x(n336), .a(n167), .b(n337) );
	nand2_5 U362 ( .x(n339), .a(n334), .b(n332) );
	nor2_5 U363 ( .x(n340), .a(n147), .b(n203) );
	aoi21_3 U364 ( .x(n344), .a(n340), .b(n345), .c(n201) );
	nor2i_5 U365 ( .x(n118), .a(n86), .b(n266) );
	nand2_2 U366 ( .x(n352), .a(n353), .b(n283) );
	nor2_5 U367 ( .x(n184), .a(n261), .b(n362) );
	oai21_5 U368 ( .x(n185), .a(n362), .b(n285), .c(n363) );
	nand2i_4 U369 ( .x(n374), .a(n329), .b(n330) );
	inv_2 U37 ( .x(n236), .a(A[19]) );
	nand2_5 U370 ( .x(n375), .a(n335), .b(n334) );
	ao21_4 U371 ( .x(n212), .a(n217), .b(n385), .c(n387) );
	nand2i_4 U372 ( .x(n395), .a(n70), .b(n270) );
	inv_5 U373 ( .x(n337), .a(n164) );
	nand2i_4 U374 ( .x(n128), .a(n406), .b(n405) );
	nand2_2 U375 ( .x(n215), .a(n372), .b(n409) );
	nand2i_4 U376 ( .x(n414), .a(n378), .b(n336) );
	inv_5 U377 ( .x(n86), .a(n267) );
	nand2i_4 U378 ( .x(n417), .a(n169), .b(n416) );
	inv_5 U379 ( .x(n378), .a(n417) );
	nor2i_0 U38 ( .x(n323), .a(B[19]), .b(n236) );
	oai21_4 U380 ( .x(n349), .a(n396), .b(n418), .c(n393) );
	nand2i_4 U381 ( .x(n415), .a(n328), .b(n379) );
	nand2i_4 U382 ( .x(n307), .a(n380), .b(n412) );
	oai21_4 U383 ( .x(n288), .a(n396), .b(n418), .c(n393) );
	inv_5 U384 ( .x(n411), .a(n295) );
	nand2i_4 U385 ( .x(n90), .a(n269), .b(n302) );
	mux2i_3 U387 ( .x(n89), .d0(n309), .sl(n407), .d1(n311) );
	mux2i_3 U388 ( .x(n79), .d0(n313), .sl(A[22]), .d1(n304) );
	nand2_3 U389 ( .x(SUM[18]), .a(n75), .b(n76) );
	nor2_3 U39 ( .x(n242), .a(n189), .b(n194) );
	nand2_3 U390 ( .x(SUM[22]), .a(n79), .b(n80) );
	nand2_3 U391 ( .x(SUM[28]), .a(n89), .b(n90) );
	exor2_5 U392 ( .x(n209), .a(B[31]), .b(n70) );
	inv_6 U393 ( .x(n162), .a(n397) );
	nand2i_4 U394 ( .x(n409), .a(n289), .b(n69) );
	nand2i_5 U395 ( .x(n82), .a(n364), .b(n69) );
	aoai211_5 U397 ( .x(n285), .a(n286), .b(n287), .c(n198), .d(n288) );
	nand2i_6 U398 ( .x(n181), .a(B[13]), .b(n251) );
	nand3i_4 U399 ( .x(n246), .a(n247), .b(n111), .c(n181) );
	nand2i_5 U400 ( .x(n342), .a(B[20]), .b(n235) );
	nand2i_4 U401 ( .x(n338), .a(n147), .b(n181) );
	nand2i_5 U402 ( .x(n263), .a(A[23]), .b(n271) );
	nand4_5 U403 ( .x(n261), .a(n262), .b(n263), .c(n264), .d(n265) );
	nand2i_6 U404 ( .x(n284), .a(n70), .b(n269) );
	nand2i_5 U405 ( .x(n381), .a(B[29]), .b(n72) );
	inv_7 U406 ( .x(n286), .a(n275) );
	nand2i_5 U407 ( .x(n389), .a(B[5]), .b(n228) );
	inv_6 U408 ( .x(n240), .a(n301) );
	inv_6 U409 ( .x(n418), .a(n419) );
	inv_2 U41 ( .x(n296), .a(n294) );
	nor2_8 U410 ( .x(n199), .a(n70), .b(B[25]) );
	or2_6 U411 ( .x(n386), .a(B[1]), .b(A[1]) );
	nand2i_8 U412 ( .x(n405), .a(n261), .b(n69) );
	exnor2_5 U413 ( .x(SUM[30]), .a(n210), .b(n65) );
	aoai211_4 U414 ( .x(n218), .a(n411), .b(n401), .c(n156), .d(n155) );
	aoai211_3 U415 ( .x(n210), .a(n285), .b(n405), .c(n355), .d(n356) );
	nand2i_5 U416 ( .x(n401), .a(n375), .b(n112) );
	nor2i_2 U417 ( .x(n313), .a(B[22]), .b(n290) );
	nand2i_2 U418 ( .x(n80), .a(n293), .b(n290) );
	inv_3 U419 ( .x(n176), .a(n386) );
	oai31_2 U42 ( .x(n295), .a(n182), .b(n165), .c(n248), .d(n296) );
	inv_0 U420 ( .x(n423), .a(n208) );
	inv_2 U421 ( .x(n424), .a(n423) );
	inv_0 U422 ( .x(n425), .a(n217) );
	inv_2 U423 ( .x(n426), .a(n425) );
	inv_0 U44 ( .x(n140), .a(n263) );
	nor2_2 U45 ( .x(n183), .a(A[22]), .b(B[22]) );
	nand2i_2 U46 ( .x(n275), .a(n183), .b(n263) );
	nand2_0 U47 ( .x(n404), .a(A[22]), .b(B[22]) );
	nand2_2 U48 ( .x(n287), .a(n404), .b(n137) );
	and3i_1 U49 ( .x(n354), .a(n352), .b(n131), .c(n124) );
	nor2i_0 U5 ( .x(n157), .a(n158), .b(n159) );
	nand2_2 U50 ( .x(n131), .a(B[26]), .b(n70) );
	nand2_0 U51 ( .x(n124), .a(B[29]), .b(n70) );
	nand2_2 U52 ( .x(n281), .a(B[27]), .b(n70) );
	nand3_1 U53 ( .x(n348), .a(n349), .b(n350), .c(n351) );
	inv_4 U54 ( .x(n350), .a(n266) );
	nand2i_2 U55 ( .x(n416), .a(B[12]), .b(n250) );
	inv_2 U56 ( .x(n363), .a(n280) );
	nand2i_0 U57 ( .x(n312), .a(B[28]), .b(n70) );
	nand2_2 U58 ( .x(n280), .a(n281), .b(n131) );
	nor2_1 U59 ( .x(n311), .a(n280), .b(n312) );
	oai21_1 U6 ( .x(n294), .a(n159), .b(n161), .c(n158) );
	inv_2 U60 ( .x(n362), .a(n310) );
	nand2_2 U61 ( .x(n310), .a(n408), .b(n72) );
	nor2_0 U62 ( .x(n322), .a(n106), .b(n103) );
	inv_2 U63 ( .x(n228), .a(A[5]) );
	inv_3 U64 ( .x(n103), .a(n318) );
	inv_2 U65 ( .x(n278), .a(n284) );
	aoi21_1 U66 ( .x(n268), .a(n347), .b(n72), .c(n278) );
	nand2i_2 U67 ( .x(n267), .a(n261), .b(n268) );
	inv_2 U68 ( .x(n197), .a(n361) );
	nand2i_2 U69 ( .x(n282), .a(n280), .b(n283) );
	exnor2_2 U7 ( .x(n302), .a(n50), .b(n49) );
	nand2_2 U70 ( .x(n359), .a(n349), .b(n351) );
	nand2i_2 U71 ( .x(n361), .a(n192), .b(n286) );
	inv_2 U72 ( .x(n360), .a(n198) );
	aoai211_1 U73 ( .x(n88), .a(n360), .b(n361), .c(n359), .d(n357) );
	nand2i_2 U74 ( .x(n127), .a(n70), .b(n260) );
	inv_2 U75 ( .x(n260), .a(B[26]) );
	nand2i_0 U76 ( .x(n319), .a(n320), .b(n321) );
	nand2_0 U77 ( .x(n99), .a(B[7]), .b(A[7]) );
	nor2i_0 U78 ( .x(n317), .a(n318), .b(n229) );
	nand2i_2 U79 ( .x(n318), .a(B[6]), .b(n230) );
	inv_2 U8 ( .x(n49), .a(n71) );
	inv_0 U80 ( .x(n230), .a(A[6]) );
	inv_2 U81 ( .x(n224), .a(B[7]) );
	inv_2 U82 ( .x(n324), .a(n229) );
	inv_4 U83 ( .x(n203), .a(n300) );
	nand2i_2 U84 ( .x(n300), .a(A[19]), .b(n144) );
	nand2i_2 U85 ( .x(n421), .a(n144), .b(n52) );
	aoi21_1 U86 ( .x(n52), .a(n219), .b(n299), .c(n297) );
	exnor2_1 U87 ( .x(n305), .a(n52), .b(n144) );
	inv_5 U88 ( .x(n144), .a(B[19]) );
	nand2i_0 U89 ( .x(n410), .a(n239), .b(n219) );
	ao21_3 U9 ( .x(n50), .a(n184), .b(n69), .c(n185) );
	nand2i_2 U90 ( .x(n376), .a(n143), .b(n377) );
	nor2i_1 U91 ( .x(n143), .a(A[19]), .b(n144) );
	nand2i_2 U92 ( .x(n377), .a(n203), .b(n297) );
	inv_0 U93 ( .x(n232), .a(B[9]) );
	nand2i_2 U94 ( .x(n402), .a(A[17]), .b(n254) );
	inv_2 U95 ( .x(n255), .a(A[16]) );
	nand2i_2 U96 ( .x(n241), .a(B[16]), .b(n255) );
	nand2i_4 U97 ( .x(n248), .a(n162), .b(n249) );
	nand2_2 U98 ( .x(n155), .a(A[16]), .b(B[16]) );
	nand2i_2 U99 ( .x(n169), .a(n60), .b(B[11]) );

endmodule


module ID_DW01_add_32_2_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire ___cell__11920_net39651, ___cell__11920_net39652, ___cell__37600_net131506,
	___cell__37600_net131507, ___cell__37600_net131508, ___cell__37600_net131509,
	___cell__37600_net131510, ___cell__37600_net131553, ___cell__37600_net131555,
	___cell__37600_net131556, ___cell__37600_net131559, ___cell__37600_net131560,
	___cell__37600_net131561, ___cell__37600_net131562, ___cell__37600_net131565,
	___cell__37600_net131566, ___cell__37600_net131568, ___cell__37600_net131570,
	___cell__37600_net131571, ___cell__37600_net131575, ___cell__37600_net131576,
	___cell__37600_net131579, ___cell__37600_net131580, ___cell__37600_net131582,
	___cell__37600_net131583, ___cell__37600_net131584, ___cell__37600_net131585,
	___cell__37600_net131586, ___cell__37600_net131596, ___cell__37600_net131608,
	___cell__37600_net131609, ___cell__37600_net131610, ___cell__37600_net131611,
	___cell__37600_net131612, ___cell__37600_net131620, ___cell__37600_net131622,
	___cell__37600_net131623, ___cell__37600_net131624, ___cell__37600_net131625,
	___cell__37600_net131627, ___cell__37600_net131630, ___cell__37600_net131631,
	___cell__37600_net131634, ___cell__37600_net131635, ___cell__37600_net131636,
	___cell__37600_net131637, ___cell__37600_net131638, ___cell__37600_net131639,
	___cell__37600_net131640, ___cell__37600_net131641, ___cell__37600_net131643,
	___cell__37600_net131645, ___cell__37600_net131652, ___cell__37600_net131672,
	___cell__37600_net131673, ___cell__37600_net131676, ___cell__37600_net131680,
	___cell__37600_net131709, ___cell__37600_net131719, ___cell__37600_net131723,
	___cell__37600_net131730, ___cell__37600_net131733, ___cell__37600_net131734,
	___cell__37600_net131735, ___cell__37600_net131736, ___cell__37600_net131737,
	___cell__37600_net131738, ___cell__37600_net131739, ___cell__37600_net131741,
	___cell__37600_net131749, ___cell__37600_net131756, ___cell__37600_net131758,
	___cell__37600_net131759, ___cell__37600_net131760, ___cell__37600_net131763,
	___cell__37600_net131766, ___cell__37600_net131767, ___cell__37600_net131770,
	___cell__37600_net131771, ___cell__37600_net131775, ___cell__37600_net131776,
	___cell__37600_net131777, ___cell__37600_net131802, ___cell__37600_net131806,
	___cell__37600_net131808, ___cell__37600_net131809, ___cell__37600_net131811,
	___cell__37600_net131819, ___cell__37600_net131821, ___cell__37600_net131823,
	___cell__37600_net131831, ___cell__37600_net131837, ___cell__37600_net131841,
	___cell__37600_net131844, ___cell__37600_net131846, ___cell__37600_net131847,
	___cell__37600_net131849, ___cell__37600_net131851, ___cell__37600_net131858,
	___cell__37600_net131859, ___cell__37600_net131861, ___cell__37600_net131866,
	___cell__37600_net131867, ___cell__37600_net131868, ___cell__37600_net131869,
	___cell__37600_net131873, n100, n101, n102, n103, n104, n105, n106, n107,
	n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
	n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
	n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
	n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
	n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
	n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
	n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
	n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
	n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
	n216, n217, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
	n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
	n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
	n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, net148303, net149302,
	net149439, net149441, net149697, net149743, net149842, net150527, net150528,
	net150977, net150978, net151157, net151423, net151639, net151640, net151781,
	net151782, net151798, net152087, net152089, net152263, net152417, net152499;


	inv_5 U10 ( .x(n183), .a(B[13]) );
	nor2i_1 U100 ( .x(n158), .a(n83), .b(n160) );
	exor2_1 U101 ( .x(SUM[14]), .a(n174), .b(n158) );
	exnor2_1 U102 ( .x(SUM[4]), .a(___cell__37600_net131624), .b(___cell__37600_net131625) );
	inv_5 U103 ( .x(n103), .a(___cell__37600_net131609) );
	nor2i_0 U104 ( .x(___cell__37600_net131611), .a(___cell__37600_net131612),
		.b(n103) );
	exor2_1 U105 ( .x(SUM[10]), .a(___cell__37600_net131608), .b(___cell__37600_net131611) );
	inv_2 U106 ( .x(___cell__37600_net131586), .a(___cell__37600_net131802) );
	nor2i_1 U107 ( .x(___cell__37600_net131575), .a(n215), .b(net152417) );
	inv_5 U108 ( .x(net152417), .a(___cell__37600_net131806) );
	exnor2_1 U109 ( .x(SUM[2]), .a(n140), .b(___cell__37600_net131584) );
	or3i_3 U11 ( .x(___cell__37600_net131756), .a(n204), .b(n137), .c(n157) );
	nor2i_1 U110 ( .x(n140), .a(n210), .b(net149842) );
	nor2i_0 U111 ( .x(___cell__37600_net131584), .a(___cell__37600_net131585),
		.b(___cell__37600_net131586) );
	exor2_1 U112 ( .x(___cell__37600_net131640), .a(net148303), .b(B[25]) );
	exnor2_1 U113 ( .x(SUM[21]), .a(n141), .b(___cell__37600_net131645) );
	aoi21_1 U114 ( .x(n141), .a(___cell__37600_net131506), .b(___cell__37600_net131507),
		.c(___cell__37600_net131508) );
	inv_0 U115 ( .x(___cell__37600_net131508), .a(___cell__37600_net131582) );
	nand2i_2 U116 ( .x(n151), .a(n187), .b(n188) );
	inv_2 U117 ( .x(n149), .a(n151) );
	exnor2_1 U118 ( .x(SUM[18]), .a(n149), .b(n171) );
	exor2_1 U119 ( .x(n169), .a(B[23]), .b(n54) );
	inv_5 U12 ( .x(n157), .a(n197) );
	inv_2 U120 ( .x(n72), .a(n52) );
	inv_4 U121 ( .x(n73), .a(B[30]) );
	inv_2 U122 ( .x(___cell__37600_net131676), .a(B[29]) );
	exnor2_1 U123 ( .x(SUM[1]), .a(n209), .b(___cell__11920_net39651) );
	nor2i_1 U124 ( .x(n209), .a(n210), .b(n208) );
	exnor2_1 U125 ( .x(SUM[5]), .a(___cell__37600_net131623), .b(___cell__37600_net131570) );
	inv_2 U126 ( .x(___cell__37600_net131623), .a(___cell__37600_net131819) );
	aoai211_1 U127 ( .x(___cell__37600_net131819), .a(___cell__37600_net131624),
		.b(n116), .c(n117), .d(n122) );
	inv_2 U128 ( .x(___cell__37600_net131624), .a(___cell__37600_net131672) );
	inv_2 U129 ( .x(n116), .a(B[4]) );
	inv_10 U13 ( .x(n163), .a(n195) );
	inv_2 U130 ( .x(n114), .a(n121) );
	inv_2 U131 ( .x(n207), .a(n175) );
	inv_2 U132 ( .x(n184), .a(B[12]) );
	exor2_1 U133 ( .x(SUM[13]), .a(n175), .b(n161) );
	inv_2 U135 ( .x(n102), .a(A[11]) );
	inv_2 U136 ( .x(n117), .a(A[4]) );
	inv_0 U137 ( .x(n185), .a(A[12]) );
	inv_10 U138 ( .x(n135), .a(B[17]) );
	oa21_2 U139 ( .x(n50), .a(___cell__37600_net131622), .b(___cell__37600_net131560),
		.c(___cell__37600_net131559) );
	inv_5 U14 ( .x(n56), .a(n90) );
	nand2_2 U140 ( .x(n51), .a(___cell__37600_net131770), .b(___cell__37600_net131771) );
	inv_5 U141 ( .x(n112), .a(B[7]) );
	inv_2 U142 ( .x(n92), .a(A[21]) );
	exor2_1 U143 ( .x(n52), .a(n74), .b(n73) );
	oai22_3 U144 ( .x(___cell__37600_net131719), .a(A[17]), .b(B[17]), .c(A[16]),
		.d(B[16]) );
	inv_2 U145 ( .x(n65), .a(A[9]) );
	exnor2_1 U146 ( .x(n53), .a(B[29]), .b(net148303) );
	inv_2 U147 ( .x(n54), .a(n126) );
	inv_2 U148 ( .x(n126), .a(A[23]) );
	aoai211_3 U149 ( .x(n55), .a(n68), .b(n67), .c(net149439), .d(___cell__37600_net131851) );
	inv_4 U15 ( .x(n49), .a(n62) );
	inv_2 U151 ( .x(n67), .a(B[28]) );
	or3i_2 U152 ( .x(n89), .a(___cell__37600_net131763), .b(net151798), .c(n57) );
	aoai211_4 U153 ( .x(___cell__37600_net131869), .a(___cell__37600_net131867),
		.b(___cell__37600_net131866), .c(net149697), .d(___cell__37600_net131766) );
	oaoi211_4 U154 ( .x(net149439), .a(net149441), .b(A[28]), .c(___cell__37600_net131637),
		.d(n51) );
	aoi21_3 U155 ( .x(net149697), .a(n56), .b(n96), .c(n98) );
	nand2i_1 U156 ( .x(n95), .a(B[21]), .b(___cell__37600_net131582) );
	or3i_5 U158 ( .x(n96), .a(___cell__37600_net131723), .b(n88), .c(n87) );
	nand2i_4 U159 ( .x(___cell__37600_net131609), .a(B[10]), .b(___cell__37600_net131709) );
	nor2_6 U16 ( .x(n62), .a(B[24]), .b(n63) );
	nor2_3 U160 ( .x(n106), .a(n103), .b(n105) );
	nand3_3 U161 ( .x(n88), .a(___cell__37600_net131758), .b(___cell__37600_net131759),
		.c(___cell__37600_net131760) );
	nand2i_4 U162 ( .x(___cell__37600_net131507), .a(A[20]), .b(n178) );
	nor2_2 U163 ( .x(n108), .a(n105), .b(___cell__37600_net131559) );
	inv_6 U164 ( .x(n105), .a(n109) );
	buf_1 U165 ( .x(n58), .a(net152263) );
	inv_5 U166 ( .x(n100), .a(n110) );
	ao31_3 U167 ( .x(n59), .a(n64), .b(n109), .c(___cell__37600_net131609),
		.d(n104) );
	exnor2_2 U169 ( .x(SUM[30]), .a(___cell__37600_net131873), .b(n72) );
	inv_6 U17 ( .x(___cell__37600_net131767), .a(n62) );
	nand4_2 U170 ( .x(n91), .a(___cell__37600_net131861), .b(___cell__37600_net131620),
		.c(___cell__37600_net131760), .d(___cell__37600_net131719) );
	inv_2 U171 ( .x(net150527), .a(___cell__37600_net131741) );
	nand2_1 U172 ( .x(n132), .a(B[1]), .b(A[1]) );
	oai211_1 U173 ( .x(n131), .a(B[1]), .b(A[1]), .c(A[0]), .d(B[0]) );
	inv_0 U174 ( .x(net151157), .a(net149439) );
	exnor2_1 U175 ( .x(n193), .a(A[12]), .b(B[12]) );
	nor2_0 U176 ( .x(n164), .a(A[12]), .b(B[12]) );
	ao21_3 U177 ( .x(net150528), .a(n108), .b(n107), .c(n101) );
	nor2_2 U178 ( .x(n107), .a(n100), .b(n103) );
	ao221_4 U179 ( .x(___cell__37600_net131637), .a(___cell__37600_net131869),
		.b(n80), .c(B[25]), .d(___cell__37600_net131869), .e(n79) );
	inv_2 U18 ( .x(n177), .a(B[27]) );
	nor2_0 U180 ( .x(n60), .a(n73), .b(n68) );
	inv_2 U181 ( .x(n61), .a(___cell__37600_net131634) );
	exor2_1 U182 ( .x(___cell__37600_net131634), .a(net148303), .b(B[28]) );
	exor2_1 U183 ( .x(SUM[6]), .a(___cell__37600_net131562), .b(n145) );
	inv_2 U184 ( .x(n63), .a(n125) );
	nor2_3 U185 ( .x(n137), .a(B[14]), .b(A[14]) );
	oai211_3 U186 ( .x(n204), .a(n163), .b(n166), .c(n162), .d(n159) );
	nand2_2 U187 ( .x(n162), .a(B[13]), .b(A[13]) );
	inv_0 U188 ( .x(n99), .a(n85) );
	nor2_3 U189 ( .x(n64), .a(n66), .b(n65) );
	nand2_1 U19 ( .x(___cell__37600_net131733), .a(A[4]), .b(B[4]) );
	inv_0 U190 ( .x(___cell__37600_net131556), .a(n64) );
	nor2i_0 U191 ( .x(n161), .a(n162), .b(n163) );
	oai21_1 U192 ( .x(n174), .a(n163), .b(n207), .c(n162) );
	nand2i_2 U193 ( .x(___cell__37600_net131596), .a(n182), .b(B[15]) );
	aoi21_3 U194 ( .x(___cell__37600_net131766), .a(n49), .b(n128), .c(n129) );
	inv_2 U195 ( .x(n68), .a(n75) );
	inv_0 U196 ( .x(___cell__37600_net131776), .a(___cell__37600_net131719) );
	exnor2_3 U197 ( .x(SUM[31]), .a(n70), .b(n69) );
	inv_2 U198 ( .x(n69), .a(net149302) );
	oaoi211_2 U199 ( .x(n70), .a(B[30]), .b(n71), .c(___cell__37600_net131873),
		.d(n60) );
	inv_2 U20 ( .x(n136), .a(n135) );
	inv_1 U200 ( .x(n71), .a(n124) );
	inv_2 U201 ( .x(net149302), .a(___cell__37600_net131627) );
	inv_0 U202 ( .x(n74), .a(net148303) );
	inv_0 U203 ( .x(n75), .a(n124) );
	inv_2 U204 ( .x(___cell__37600_net131851), .a(n76) );
	inv_0 U205 ( .x(n77), .a(net148303) );
	exor2_1 U206 ( .x(SUM[23]), .a(___cell__37600_net131643), .b(n169) );
	nor2i_0 U207 ( .x(n144), .a(___cell__37600_net131559), .b(___cell__37600_net131560) );
	oai211_2 U208 ( .x(___cell__37600_net131808), .a(___cell__37600_net131735),
		.b(___cell__37600_net131734), .c(___cell__37600_net131809), .d(___cell__37600_net131739) );
	oai211_2 U209 ( .x(___cell__37600_net131735), .a(___cell__37600_net131630),
		.b(___cell__37600_net131736), .c(___cell__37600_net131737), .d(___cell__37600_net131738) );
	nand2_2 U21 ( .x(___cell__37600_net131758), .a(A[17]), .b(n136) );
	inv_2 U210 ( .x(n80), .a(n124) );
	inv_0 U211 ( .x(___cell__37600_net131639), .a(___cell__37600_net131869) );
	nand2_1 U212 ( .x(___cell__37600_net131846), .a(B[25]), .b(net148303) );
	inv_0 U213 ( .x(n124), .a(A[31]) );
	inv_0 U214 ( .x(n81), .a(___cell__37600_net131847) );
	nand2_5 U215 ( .x(___cell__37600_net131760), .a(A[18]), .b(n139) );
	inv_3 U216 ( .x(n138), .a(B[18]) );
	nand2i_4 U217 ( .x(n188), .a(___cell__37600_net131719), .b(n154) );
	inv_0 U218 ( .x(n201), .a(n203) );
	nand2_0 U219 ( .x(___cell__37600_net131837), .a(A[18]), .b(n139) );
	nand2i_2 U22 ( .x(___cell__37600_net131861), .a(n181), .b(n203) );
	aoi21_1 U220 ( .x(___cell__37600_net131509), .a(___cell__37600_net131510),
		.b(___cell__37600_net131506), .c(n213) );
	nor2i_1 U221 ( .x(n156), .a(___cell__37600_net131596), .b(n157) );
	nor2_0 U222 ( .x(___cell__37600_net131510), .a(___cell__37600_net131583),
		.b(net151798) );
	inv_0 U223 ( .x(n82), .a(n159) );
	inv_2 U224 ( .x(n83), .a(n82) );
	inv_0 U225 ( .x(___cell__37600_net131643), .a(net149697) );
	inv_0 U226 ( .x(___cell__37600_net131580), .a(___cell__37600_net131763) );
	nand2_5 U227 ( .x(n87), .a(___cell__37600_net131756), .b(n86) );
	and2_3 U228 ( .x(n86), .a(___cell__37600_net131620), .b(___cell__37600_net131596) );
	nor2i_3 U229 ( .x(n84), .a(___cell__37600_net131620), .b(net152263) );
	oa22_3 U23 ( .x(net152263), .a(B[18]), .b(A[18]), .c(B[19]), .d(A[19]) );
	nand2_1 U230 ( .x(n94), .a(___cell__37600_net131582), .b(n92) );
	inv_2 U231 ( .x(n97), .a(n93) );
	exor2_1 U232 ( .x(___cell__37600_net131645), .a(A[21]), .b(n97) );
	inv_0 U233 ( .x(n85), .a(A[22]) );
	nand2_1 U234 ( .x(___cell__37600_net131579), .a(A[22]), .b(B[22]) );
	ao211_5 U235 ( .x(___cell__37600_net131831), .a(net150527), .b(___cell__37600_net131808),
		.c(net150528), .d(n59) );
	nand2i_4 U236 ( .x(___cell__37600_net131723), .a(___cell__37600_net131749),
		.b(___cell__37600_net131831) );
	inv_0 U237 ( .x(___cell__37600_net131730), .a(___cell__37600_net131831) );
	and3i_2 U238 ( .x(n104), .a(n105), .b(n78), .c(A[10]) );
	inv_0 U239 ( .x(n111), .a(n102) );
	nand2_2 U24 ( .x(___cell__37600_net131582), .a(A[20]), .b(B[20]) );
	exor2_1 U240 ( .x(___cell__37600_net131652), .a(B[11]), .b(n111) );
	or3i_2 U241 ( .x(___cell__37600_net131741), .a(n106), .b(n100), .c(___cell__37600_net131560) );
	oai21_1 U242 ( .x(___cell__37600_net131608), .a(n50), .b(n100), .c(___cell__37600_net131556) );
	nor2i_0 U243 ( .x(___cell__37600_net131555), .a(___cell__37600_net131556),
		.b(n100) );
	inv_0 U244 ( .x(___cell__37600_net131622), .a(___cell__37600_net131808) );
	aoi21_3 U245 ( .x(___cell__37600_net131739), .a(n119), .b(n120), .c(___cell__37600_net131553) );
	nor2i_1 U246 ( .x(___cell__37600_net131553), .a(A[7]), .b(n112) );
	nand2i_6 U247 ( .x(___cell__37600_net131738), .a(A[7]), .b(n112) );
	aoi21_2 U248 ( .x(n120), .a(___cell__37600_net131571), .b(___cell__37600_net131733),
		.c(n115) );
	nor2_1 U249 ( .x(n115), .a(B[5]), .b(A[5]) );
	nand2i_2 U25 ( .x(n196), .a(A[12]), .b(n184) );
	nor2_8 U250 ( .x(n119), .a(___cell__37600_net131566), .b(net152087) );
	aoi21_1 U251 ( .x(___cell__37600_net131565), .a(n217), .b(B[7]), .c(___cell__37600_net131566) );
	nand2i_4 U252 ( .x(___cell__37600_net131734), .a(n114), .b(n113) );
	oai21_1 U253 ( .x(___cell__37600_net131562), .a(n114), .b(___cell__37600_net131623),
		.c(___cell__37600_net131571) );
	nor2i_0 U254 ( .x(___cell__37600_net131570), .a(___cell__37600_net131571),
		.b(n114) );
	aoi21_4 U255 ( .x(___cell__37600_net131737), .a(n116), .b(n117), .c(net152417) );
	aoai211_4 U256 ( .x(___cell__37600_net131873), .a(n123), .b(___cell__37600_net131676),
		.c(___cell__37600_net131631), .d(___cell__37600_net131859) );
	inv_2 U257 ( .x(n123), .a(A[31]) );
	aoai211_1 U259 ( .x(___cell__37600_net131635), .a(___cell__37600_net131680),
		.b(n124), .c(___cell__37600_net131847), .d(___cell__37600_net131770) );
	nand2_1 U26 ( .x(___cell__37600_net131770), .a(B[26]), .b(net148303) );
	inv_5 U260 ( .x(net149441), .a(___cell__37600_net131868) );
	nand2i_4 U261 ( .x(___cell__37600_net131868), .a(___cell__37600_net131680),
		.b(___cell__37600_net131849) );
	inv_0 U262 ( .x(___cell__37600_net131847), .a(___cell__37600_net131637) );
	exor2_1 U263 ( .x(SUM[26]), .a(n81), .b(___cell__37600_net131638) );
	nand2_3 U264 ( .x(___cell__37600_net131636), .a(___cell__37600_net131771),
		.b(___cell__37600_net131849) );
	exor2_2 U265 ( .x(___cell__37600_net131627), .a(net148303), .b(B[31]) );
	nor2i_6 U266 ( .x(n128), .a(A[23]), .b(n127) );
	inv_10 U267 ( .x(n127), .a(B[23]) );
	nand2i_4 U268 ( .x(___cell__37600_net131866), .a(n127), .b(___cell__37600_net131767) );
	nand2i_4 U269 ( .x(___cell__37600_net131867), .a(n126), .b(___cell__37600_net131767) );
	nand2_2 U27 ( .x(___cell__37600_net131771), .a(B[27]), .b(net148303) );
	inv_0 U270 ( .x(___cell__37600_net131821), .a(___cell__37600_net131767) );
	inv_0 U271 ( .x(n125), .a(A[24]) );
	nand2_2 U272 ( .x(___cell__37600_net131844), .a(A[24]), .b(B[24]) );
	inv_0 U273 ( .x(___cell__37600_net131673), .a(___cell__37600_net131630) );
	nand2_2 U274 ( .x(___cell__37600_net131585), .a(A[2]), .b(B[2]) );
	inv_0 U275 ( .x(net150977), .a(A[1]) );
	inv_0 U276 ( .x(net151639), .a(A[0]) );
	nand2_0 U277 ( .x(___cell__11920_net39651), .a(net151640), .b(B[0]) );
	nor2_0 U278 ( .x(___cell__11920_net39652), .a(B[0]), .b(net151640) );
	oa211_1 U279 ( .x(net149842), .a(B[1]), .b(net150978), .c(net151640), .d(B[0]) );
	nor2i_1 U28 ( .x(n76), .a(B[28]), .b(n77) );
	nand2i_4 U280 ( .x(___cell__37600_net131806), .a(B[3]), .b(n133) );
	exor2_1 U281 ( .x(___cell__37600_net131625), .a(A[4]), .b(B[4]) );
	oai21_1 U282 ( .x(___cell__37600_net131672), .a(___cell__37600_net131673),
		.b(net152417), .c(n215) );
	exnor2_1 U283 ( .x(SUM[25]), .a(___cell__37600_net131639), .b(___cell__37600_net131640) );
	exnor2_1 U284 ( .x(SUM[8]), .a(___cell__37600_net131622), .b(n144) );
	and2_2 U285 ( .x(net152499), .a(A[6]), .b(B[6]) );
	inv_0 U286 ( .x(___cell__37600_net131568), .a(net152499) );
	mux2i_1 U287 ( .x(SUM[12]), .d0(n165), .sl(___cell__37600_net131730), .d1(n193) );
	aoai211_1 U288 ( .x(n175), .a(n185), .b(n184), .c(___cell__37600_net131730),
		.d(n166) );
	inv_6 U289 ( .x(___cell__37600_net131709), .a(A[10]) );
	inv_2 U29 ( .x(net148303), .a(n123) );
	nand3_0 U290 ( .x(n199), .a(___cell__37600_net131758), .b(___cell__37600_net131759),
		.c(___cell__37600_net131760) );
	buf_3 U291 ( .x(n134), .a(B[8]) );
	exor2_1 U292 ( .x(SUM[3]), .a(___cell__37600_net131630), .b(___cell__37600_net131575) );
	inv_2 U293 ( .x(n182), .a(A[15]) );
	inv_0 U294 ( .x(net151781), .a(___cell__37600_net131723) );
	aoi21_1 U296 ( .x(n152), .a(n153), .b(n154), .c(n155) );
	oai22_1 U297 ( .x(n187), .a(n135), .b(n186), .c(n201), .d(n211) );
	nand2i_0 U298 ( .x(n143), .a(n186), .b(n154) );
	inv_0 U299 ( .x(___cell__37600_net131841), .a(___cell__37600_net131620) );
	nand2i_2 U30 ( .x(___cell__37600_net131809), .a(___cell__37600_net131566),
		.b(net152499) );
	nand2_1 U300 ( .x(___cell__37600_net131759), .a(A[16]), .b(B[16]) );
	nand2_0 U301 ( .x(n186), .a(A[16]), .b(B[16]) );
	inv_2 U303 ( .x(net151640), .a(net151639) );
	or3i_1 U305 ( .x(n206), .a(net151782), .b(n198), .c(n199) );
	inv_0 U306 ( .x(net151423), .a(___cell__37600_net131643) );
	exor2_1 U307 ( .x(n170), .a(B[19]), .b(A[19]) );
	inv_2 U308 ( .x(net150978), .a(net150977) );
	exnor2_1 U309 ( .x(n189), .a(A[9]), .b(net149743) );
	nand2i_2 U31 ( .x(n121), .a(B[5]), .b(n118) );
	inv_4 U310 ( .x(n139), .a(n138) );
	nand2_0 U311 ( .x(n198), .a(___cell__37600_net131756), .b(___cell__37600_net131596) );
	nand2_2 U312 ( .x(___cell__37600_net131571), .a(A[5]), .b(B[5]) );
	inv_0 U313 ( .x(n179), .a(B[16]) );
	nand2i_0 U314 ( .x(n153), .a(B[16]), .b(n180) );
	ao21_3 U315 ( .x(n203), .a(A[16]), .b(B[16]), .c(B[17]) );
	inv_0 U316 ( .x(n160), .a(n194) );
	nand2_0 U317 ( .x(___cell__37600_net131612), .a(A[10]), .b(n78) );
	mux2i_1 U318 ( .x(SUM[7]), .d0(___cell__37600_net131565), .sl(___cell__37600_net131561),
		.d1(n190) );
	exnor2_1 U319 ( .x(n190), .a(n217), .b(B[7]) );
	nand2_1 U32 ( .x(___cell__37600_net131576), .a(A[3]), .b(B[3]) );
	oai31_1 U320 ( .x(n200), .a(___cell__37600_net131775), .b(___cell__37600_net131776),
		.c(___cell__37600_net131777), .d(n58) );
	nand2_0 U321 ( .x(n210), .a(net150978), .b(B[1]) );
	nor2_0 U322 ( .x(n208), .a(B[1]), .b(net150978) );
	nor2i_3 U323 ( .x(n148), .a(n139), .b(n149) );
	exor2_1 U324 ( .x(n171), .a(A[18]), .b(n139) );
	oaoi211_1 U325 ( .x(n150), .a(n139), .b(n151), .c(A[18]), .d(n148) );
	nand4_1 U326 ( .x(___cell__37600_net131749), .a(n197), .b(n195), .c(n196),
		.d(n194) );
	nand2i_6 U327 ( .x(___cell__37600_net131849), .a(net148303), .b(n177) );
	nand2i_2 U328 ( .x(n154), .a(n198), .b(net151782) );
	inv_2 U329 ( .x(net151782), .a(net151781) );
	inv_7 U33 ( .x(___cell__37600_net131566), .a(___cell__37600_net131738) );
	inv_4 U330 ( .x(___cell__37600_net131631), .a(n55) );
	exnor2_1 U331 ( .x(SUM[29]), .a(n55), .b(n53) );
	inv_0 U332 ( .x(n211), .a(A[17]) );
	inv_2 U333 ( .x(n181), .a(A[17]) );
	exnor2_3 U334 ( .x(SUM[19]), .a(n150), .b(n170) );
	inv_0 U335 ( .x(n212), .a(net152089) );
	inv_2 U336 ( .x(n213), .a(n212) );
	oa211_4 U337 ( .x(net152089), .a(A[21]), .b(n97), .c(n94), .d(n95) );
	aoai211_2 U338 ( .x(___cell__37600_net131630), .a(n131), .b(n132), .c(___cell__37600_net131586),
		.d(___cell__37600_net131585) );
	inv_0 U339 ( .x(n214), .a(___cell__37600_net131576) );
	buf_2 U34 ( .x(net149743), .a(B[9]) );
	inv_2 U340 ( .x(n215), .a(n214) );
	nand2_3 U341 ( .x(___cell__37600_net131620), .a(A[19]), .b(B[19]) );
	inv_0 U342 ( .x(n216), .a(A[7]) );
	inv_2 U343 ( .x(n217), .a(n216) );
	buf_2 U35 ( .x(n78), .a(B[10]) );
	nor2i_0 U36 ( .x(n101), .a(B[11]), .b(n102) );
	nor2i_0 U37 ( .x(n192), .a(n179), .b(n154) );
	exnor2_1 U38 ( .x(n191), .a(n154), .b(n179) );
	inv_2 U40 ( .x(___cell__37600_net131777), .a(___cell__37600_net131837) );
	inv_0 U41 ( .x(___cell__37600_net131775), .a(___cell__37600_net131861) );
	nand2i_2 U42 ( .x(n205), .a(n200), .b(n206) );
	inv_2 U43 ( .x(n176), .a(A[8]) );
	nand2i_2 U44 ( .x(___cell__37600_net131811), .a(B[8]), .b(n176) );
	nand2_2 U45 ( .x(___cell__37600_net131559), .a(A[8]), .b(n134) );
	inv_2 U46 ( .x(n180), .a(A[16]) );
	nand2_2 U47 ( .x(___cell__37600_net131858), .a(B[23]), .b(n54) );
	nand2i_4 U48 ( .x(n197), .a(B[15]), .b(n182) );
	inv_4 U49 ( .x(n113), .a(net152087) );
	oa21_3 U5 ( .x(n98), .a(net152089), .b(___cell__37600_net131823), .c(___cell__37600_net131763) );
	nor2_6 U50 ( .x(net152087), .a(B[6]), .b(A[6]) );
	nand2_2 U51 ( .x(n159), .a(A[14]), .b(B[14]) );
	inv_2 U52 ( .x(n66), .a(net149743) );
	nand2i_2 U53 ( .x(n110), .a(B[9]), .b(n65) );
	inv_2 U54 ( .x(n133), .a(A[3]) );
	inv_2 U55 ( .x(___cell__37600_net131736), .a(___cell__37600_net131576) );
	inv_4 U56 ( .x(n130), .a(A[2]) );
	nand2i_2 U57 ( .x(___cell__37600_net131802), .a(B[2]), .b(n130) );
	inv_2 U58 ( .x(n129), .a(___cell__37600_net131844) );
	inv_5 U59 ( .x(n178), .a(B[20]) );
	or2_6 U6 ( .x(___cell__37600_net131763), .a(B[22]), .b(n99) );
	or3i_2 U60 ( .x(n90), .a(n91), .b(n84), .c(n89) );
	inv_2 U61 ( .x(n57), .a(___cell__37600_net131507) );
	inv_2 U62 ( .x(___cell__37600_net131823), .a(___cell__37600_net131579) );
	inv_3 U63 ( .x(n93), .a(B[21]) );
	nand2_2 U64 ( .x(___cell__37600_net131859), .a(B[29]), .b(net148303) );
	inv_2 U65 ( .x(n118), .a(A[5]) );
	nand2i_2 U66 ( .x(n122), .a(n116), .b(___cell__37600_net131672) );
	nand2_2 U67 ( .x(n166), .a(A[12]), .b(B[12]) );
	inv_5 U68 ( .x(___cell__37600_net131680), .a(B[26]) );
	exnor2_1 U69 ( .x(SUM[27]), .a(___cell__37600_net131635), .b(___cell__37600_net131636) );
	nand2i_4 U7 ( .x(n109), .a(B[11]), .b(n102) );
	exnor2_1 U70 ( .x(SUM[28]), .a(net151157), .b(n61) );
	aoi21_1 U71 ( .x(___cell__37600_net131561), .a(___cell__37600_net131562),
		.b(n113), .c(net152499) );
	inv_2 U72 ( .x(n79), .a(___cell__37600_net131846) );
	exor2_1 U73 ( .x(___cell__37600_net131638), .a(net148303), .b(B[26]) );
	nor2i_1 U74 ( .x(n165), .a(n166), .b(n164) );
	mux2i_1 U75 ( .x(n142), .d0(n191), .sl(A[16]), .d1(n192) );
	nand2_2 U76 ( .x(SUM[16]), .a(n142), .b(n143) );
	exor2_1 U77 ( .x(SUM[20]), .a(___cell__37600_net131506), .b(n147) );
	nand2i_2 U78 ( .x(___cell__37600_net131506), .a(___cell__37600_net131841),
		.b(n205) );
	nor2i_1 U79 ( .x(n147), .a(___cell__37600_net131582), .b(___cell__37600_net131583) );
	and2_3 U8 ( .x(net151798), .a(n92), .b(n93) );
	inv_2 U80 ( .x(___cell__37600_net131583), .a(___cell__37600_net131507) );
	inv_2 U81 ( .x(___cell__37600_net131560), .a(___cell__37600_net131811) );
	mux2i_1 U82 ( .x(SUM[9]), .d0(___cell__37600_net131555), .sl(n50), .d1(n189) );
	exor2_1 U83 ( .x(n172), .a(A[17]), .b(n136) );
	inv_2 U84 ( .x(n155), .a(n186) );
	exnor2_1 U85 ( .x(SUM[17]), .a(n152), .b(n172) );
	nor2i_1 U86 ( .x(SUM[0]), .a(___cell__11920_net39651), .b(___cell__11920_net39652) );
	exnor2_1 U87 ( .x(SUM[11]), .a(n167), .b(___cell__37600_net131652) );
	aoi21_1 U88 ( .x(n167), .a(___cell__37600_net131608), .b(___cell__37600_net131609),
		.c(___cell__37600_net131610) );
	inv_2 U89 ( .x(___cell__37600_net131610), .a(___cell__37600_net131612) );
	nand2i_3 U9 ( .x(n195), .a(A[13]), .b(n183) );
	exnor2_1 U90 ( .x(SUM[22]), .a(___cell__37600_net131509), .b(n146) );
	nor2i_1 U91 ( .x(n146), .a(___cell__37600_net131579), .b(___cell__37600_net131580) );
	nand2i_0 U92 ( .x(n168), .a(___cell__37600_net131821), .b(___cell__37600_net131844) );
	aoai211_1 U93 ( .x(___cell__37600_net131641), .a(n126), .b(n127), .c(net151423),
		.d(___cell__37600_net131858) );
	exnor2_1 U94 ( .x(SUM[24]), .a(___cell__37600_net131641), .b(n168) );
	exor2_1 U95 ( .x(SUM[15]), .a(n173), .b(n156) );
	oai21_1 U96 ( .x(n173), .a(n160), .b(n202), .c(n83) );
	inv_2 U97 ( .x(n194), .a(n137) );
	nor2i_0 U98 ( .x(n145), .a(___cell__37600_net131568), .b(net152087) );
	inv_2 U99 ( .x(n202), .a(n174) );

endmodule


module ID_DW01_add_32_1_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
	n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
	n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
	n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
	n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
	n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
	n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
	n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
	n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
	n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
	n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
	n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
	n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
	n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
	n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339,
	n340, n341, n342, n343, n344, n345, n346, n347, n49, n50, n51, n52, n53,
	n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
	n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
	n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
	n96, n97, n98, n99;


	ao21_3 U10 ( .x(n277), .a(n217), .b(n218), .c(n106) );
	nand2i_2 U100 ( .x(n173), .a(B[30]), .b(n170) );
	nor2i_1 U101 ( .x(n177), .a(n178), .b(n176) );
	ao21_1 U102 ( .x(n191), .a(n314), .b(n79), .c(n316) );
	inv_2 U103 ( .x(n219), .a(A[4]) );
	inv_2 U104 ( .x(n316), .a(n105) );
	nand2_2 U105 ( .x(n105), .a(A[4]), .b(B[4]) );
	inv_2 U106 ( .x(n321), .a(n191) );
	inv_2 U107 ( .x(n106), .a(n314) );
	inv_5 U108 ( .x(n62), .a(B[13]) );
	nand2_0 U109 ( .x(n110), .a(n302), .b(n146) );
	nand2i_3 U11 ( .x(n308), .a(B[6]), .b(n216) );
	nand2i_2 U110 ( .x(n302), .a(n149), .b(n325) );
	nand2i_0 U111 ( .x(n301), .a(n282), .b(n283) );
	inv_2 U112 ( .x(n282), .a(n152) );
	inv_2 U113 ( .x(n322), .a(n127) );
	exnor2_3 U114 ( .x(SUM[27]), .a(n199), .b(n53) );
	exor2_1 U115 ( .x(SUM[7]), .a(n188), .b(n189) );
	ao21_1 U116 ( .x(n188), .a(n190), .b(n66), .c(n55) );
	exnor2_1 U117 ( .x(SUM[8]), .a(n186), .b(n187) );
	nand2i_2 U118 ( .x(n187), .a(n230), .b(n232) );
	exor2_1 U119 ( .x(SUM[12]), .a(n212), .b(n145) );
	nor2i_3 U12 ( .x(n157), .a(B[7]), .b(n158) );
	oai21_1 U120 ( .x(n212), .a(n305), .b(n150), .c(n85) );
	inv_2 U121 ( .x(n305), .a(n109) );
	inv_0 U122 ( .x(n150), .a(n226) );
	nor2i_0 U123 ( .x(n145), .a(n146), .b(n147) );
	inv_0 U124 ( .x(n147), .a(n325) );
	inv_2 U125 ( .x(n265), .a(n139) );
	nor2i_1 U126 ( .x(n135), .a(n136), .b(n137) );
	inv_2 U127 ( .x(n137), .a(n337) );
	exor2_1 U128 ( .x(n210), .a(B[19]), .b(n87) );
	nand2_2 U129 ( .x(n209), .a(n328), .b(n336) );
	inv_0 U13 ( .x(n239), .a(B[18]) );
	exor2_1 U130 ( .x(SUM[19]), .a(n209), .b(n210) );
	exor2_1 U131 ( .x(n207), .a(B[20]), .b(n88) );
	inv_2 U132 ( .x(n240), .a(B[19]) );
	inv_2 U133 ( .x(n328), .a(n267) );
	oai22_1 U134 ( .x(n206), .a(n328), .b(n240), .c(n117), .d(n170) );
	exor2_1 U136 ( .x(SUM[9]), .a(n185), .b(n98) );
	oai21_1 U137 ( .x(n185), .a(n320), .b(n230), .c(n232) );
	inv_2 U138 ( .x(n230), .a(n319) );
	nor2i_0 U139 ( .x(n98), .a(n99), .b(n100) );
	nand2_2 U14 ( .x(n245), .a(B[18]), .b(n88) );
	inv_5 U140 ( .x(n100), .a(n231) );
	exor2_1 U141 ( .x(SUM[17]), .a(n211), .b(n132) );
	nor2i_1 U142 ( .x(SUM[0]), .a(n89), .b(n90) );
	exor2_1 U143 ( .x(SUM[11]), .a(n109), .b(n148) );
	nand2_2 U144 ( .x(SUM[22]), .a(n96), .b(n97) );
	nand2i_2 U146 ( .x(n97), .a(n263), .b(n261) );
	exnor2_1 U147 ( .x(SUM[15]), .a(n114), .b(n138) );
	aoi21_1 U148 ( .x(n114), .a(n115), .b(n109), .c(n116) );
	nor2i_1 U149 ( .x(n138), .a(n139), .b(n140) );
	inv_2 U15 ( .x(n163), .a(B[13]) );
	inv_5 U150 ( .x(n140), .a(n327) );
	exor2_1 U151 ( .x(SUM[6]), .a(n190), .b(n101) );
	exnor2_1 U152 ( .x(SUM[14]), .a(n111), .b(n141) );
	exor2_1 U153 ( .x(SUM[4]), .a(n79), .b(n104) );
	nor2i_0 U154 ( .x(n104), .a(n105), .b(n106) );
	exor2_1 U155 ( .x(SUM[10]), .a(n213), .b(n151) );
	oai21_1 U156 ( .x(n213), .a(n320), .b(n229), .c(n51) );
	inv_2 U157 ( .x(n320), .a(n186) );
	nor2i_0 U158 ( .x(n151), .a(n152), .b(n153) );
	exor2_1 U159 ( .x(SUM[3]), .a(n74), .b(n123) );
	nor2i_1 U16 ( .x(n162), .a(A[13]), .b(n163) );
	inv_2 U160 ( .x(n313), .a(n130) );
	nor2i_1 U161 ( .x(n123), .a(n124), .b(n125) );
	inv_2 U162 ( .x(n131), .a(n311) );
	nor2i_1 U163 ( .x(n129), .a(n130), .b(n131) );
	exor2_1 U164 ( .x(SUM[2]), .a(n80), .b(n129) );
	inv_2 U165 ( .x(n323), .a(n250) );
	nand2i_2 U166 ( .x(n202), .a(n323), .b(n254) );
	mux2i_1 U167 ( .x(n94), .d0(n275), .sl(B[21]), .d1(n169) );
	inv_0 U169 ( .x(n93), .a(n345) );
	nor2_1 U17 ( .x(n278), .a(B[22]), .b(B[21]) );
	nand2_2 U170 ( .x(SUM[18]), .a(n91), .b(n92) );
	nand3i_1 U171 ( .x(n92), .a(n347), .b(n87), .c(n338) );
	inv_2 U172 ( .x(n338), .a(n269) );
	nand3i_1 U173 ( .x(n204), .a(n307), .b(n346), .c(n262) );
	inv_2 U174 ( .x(n307), .a(n263) );
	inv_3 U176 ( .x(n70), .a(n59) );
	nor2i_1 U177 ( .x(n154), .a(n57), .b(n156) );
	exnor2_1 U178 ( .x(SUM[1]), .a(n154), .b(n89) );
	inv_2 U179 ( .x(n108), .a(n225) );
	nand2i_3 U18 ( .x(n258), .a(n289), .b(n268) );
	aoi21_1 U180 ( .x(n107), .a(n108), .b(n109), .c(n110) );
	inv_0 U181 ( .x(n58), .a(A[14]) );
	oa21_1 U183 ( .x(n51), .a(n100), .b(n232), .c(n99) );
	exnor2_1 U184 ( .x(n53), .a(B[27]), .b(n87) );
	aoai211_4 U185 ( .x(n171), .a(n75), .b(n256), .c(n258), .d(n259) );
	exnor2_1 U187 ( .x(n54), .a(B[28]), .b(n87) );
	aoi22_2 U188 ( .x(n172), .a(B[30]), .b(n88), .c(n174), .d(n173) );
	nand2i_2 U189 ( .x(n109), .a(n301), .b(n304) );
	nand2_2 U19 ( .x(n289), .a(B[20]), .b(B[19]) );
	aoai211_3 U190 ( .x(n304), .a(n343), .b(n317), .c(n342), .d(n279) );
	oai21_1 U191 ( .x(SUM[21]), .a(n93), .b(n94), .c(n95) );
	inv_5 U192 ( .x(n69), .a(A[3]) );
	nor2i_2 U193 ( .x(n183), .a(B[21]), .b(n184) );
	nand3i_5 U194 ( .x(n306), .a(B[21]), .b(n184), .c(n345) );
	nand2_1 U195 ( .x(n152), .a(A[10]), .b(B[10]) );
	nor2i_3 U196 ( .x(n67), .a(n68), .b(A[1]) );
	oai21_3 U197 ( .x(n271), .a(n100), .b(n232), .c(n99) );
	inv_0 U198 ( .x(n56), .a(n218) );
	nand2i_0 U199 ( .x(n337), .a(B[16]), .b(n170) );
	or3i_2 U20 ( .x(n249), .a(n250), .b(n248), .c(n247) );
	nand2_0 U200 ( .x(n136), .a(B[16]), .b(n87) );
	buf_1 U201 ( .x(n57), .a(n155) );
	nor2_1 U202 ( .x(n175), .a(B[5]), .b(A[5]) );
	and2_5 U203 ( .x(n143), .a(n58), .b(n237) );
	and2_5 U204 ( .x(n256), .a(n288), .b(n287) );
	nand2i_2 U205 ( .x(n66), .a(B[6]), .b(n216) );
	inv_2 U206 ( .x(n72), .a(B[0]) );
	nor2i_5 U207 ( .x(n60), .a(n62), .b(n61) );
	inv_0 U208 ( .x(n159), .a(n60) );
	inv_2 U209 ( .x(n61), .a(n236) );
	nor2i_2 U21 ( .x(n279), .a(n280), .b(n229) );
	inv_0 U210 ( .x(n236), .a(A[13]) );
	or3i_2 U211 ( .x(n63), .a(n257), .b(n265), .c(n266) );
	or3i_3 U212 ( .x(n119), .a(n257), .b(n265), .c(n266) );
	inv_7 U213 ( .x(n342), .a(n341) );
	ao211_5 U214 ( .x(n75), .a(n304), .b(n81), .c(n233), .d(n140) );
	or3i_4 U215 ( .x(n330), .a(n82), .b(n222), .c(n293) );
	nor2_2 U216 ( .x(n76), .a(n69), .b(n77) );
	inv_0 U217 ( .x(n64), .a(B[13]) );
	inv_2 U218 ( .x(n65), .a(n64) );
	nand2i_0 U219 ( .x(n186), .a(n179), .b(n341) );
	nand2_2 U22 ( .x(n343), .a(n180), .b(n181) );
	nand2_2 U220 ( .x(n310), .a(n77), .b(n69) );
	exnor2_3 U221 ( .x(SUM[28]), .a(n198), .b(n54) );
	inv_3 U222 ( .x(n312), .a(n67) );
	inv_0 U223 ( .x(n89), .a(n70) );
	nor2i_0 U224 ( .x(n141), .a(n142), .b(n143) );
	oai31_1 U225 ( .x(n116), .a(n160), .b(n143), .c(n60), .d(n142) );
	nand2_5 U226 ( .x(n329), .a(n250), .b(n201) );
	nand4i_3 U227 ( .x(n174), .a(n161), .b(n330), .c(n331), .d(n332) );
	buf_4 U228 ( .x(n71), .a(B[12]) );
	nand2i_2 U229 ( .x(n333), .a(n295), .b(n82) );
	nand2_2 U23 ( .x(n283), .a(n271), .b(n280) );
	exnor2_1 U230 ( .x(SUM[25]), .a(n82), .b(n202) );
	inv_3 U231 ( .x(n83), .a(n184) );
	oai211_4 U232 ( .x(n201), .a(n184), .b(n120), .c(n290), .d(n345) );
	inv_2 U233 ( .x(n77), .a(B[3]) );
	exor2_1 U234 ( .x(n189), .a(B[7]), .b(A[7]) );
	inv_2 U235 ( .x(n158), .a(A[7]) );
	inv_0 U236 ( .x(n73), .a(n195) );
	inv_2 U237 ( .x(n74), .a(n73) );
	nand2_5 U238 ( .x(n232), .a(A[8]), .b(B[8]) );
	inv_4 U239 ( .x(n220), .a(A[8]) );
	nand2i_2 U24 ( .x(n280), .a(B[10]), .b(n228) );
	nor2i_1 U240 ( .x(n117), .a(n118), .b(n63) );
	exor2_1 U241 ( .x(SUM[16]), .a(n63), .b(n135) );
	nand2i_0 U242 ( .x(n336), .a(n170), .b(n63) );
	ao21_3 U243 ( .x(n211), .a(n337), .b(n63), .c(n324) );
	inv_0 U244 ( .x(n156), .a(n312) );
	ao211_3 U245 ( .x(n257), .a(n304), .b(n81), .c(n140), .d(n233) );
	nand2_2 U246 ( .x(n253), .a(B[27]), .b(n88) );
	inv_0 U247 ( .x(n124), .a(n76) );
	ao21_4 U248 ( .x(n192), .a(n310), .b(n195), .c(n76) );
	inv_0 U249 ( .x(n125), .a(n310) );
	inv_0 U25 ( .x(n228), .a(A[10]) );
	nand2_1 U250 ( .x(n318), .a(B[5]), .b(A[5]) );
	nand2_0 U251 ( .x(n178), .a(n56), .b(A[5]) );
	nor2_0 U252 ( .x(n176), .a(n56), .b(A[5]) );
	nand2i_2 U253 ( .x(n334), .a(n50), .b(n170) );
	inv_2 U254 ( .x(n248), .a(B[26]) );
	nor2_1 U255 ( .x(n164), .a(B[13]), .b(A[13]) );
	aoi21_1 U256 ( .x(n144), .a(A[13]), .b(n65), .c(n60) );
	inv_0 U257 ( .x(n78), .a(n192) );
	inv_2 U258 ( .x(n79), .a(n78) );
	nand2_3 U259 ( .x(n99), .a(A[9]), .b(B[9]) );
	inv_2 U26 ( .x(n128), .a(n334) );
	oai21_1 U260 ( .x(n80), .a(n156), .b(n89), .c(n57) );
	inv_4 U261 ( .x(n216), .a(A[6]) );
	inv_2 U262 ( .x(n235), .a(A[11]) );
	nand2_1 U263 ( .x(n149), .a(A[11]), .b(B[11]) );
	inv_0 U264 ( .x(n115), .a(n233) );
	nand2i_6 U265 ( .x(n327), .a(n86), .b(n224) );
	nand2i_2 U266 ( .x(n281), .a(n282), .b(n283) );
	oai211_1 U267 ( .x(n95), .a(n93), .b(n83), .c(n88), .d(B[21]) );
	nand2_1 U268 ( .x(n346), .a(n309), .b(n83) );
	aoi21_1 U269 ( .x(n167), .a(n298), .b(n83), .c(n299) );
	inv_2 U27 ( .x(n247), .a(B[27]) );
	oai211_4 U270 ( .x(n82), .a(n184), .b(n120), .c(n290), .d(n345) );
	nand2i_2 U271 ( .x(n311), .a(A[2]), .b(n214) );
	nand2_2 U272 ( .x(n130), .a(B[2]), .b(A[2]) );
	inv_0 U273 ( .x(n84), .a(n149) );
	inv_2 U274 ( .x(n85), .a(n84) );
	nor2_0 U275 ( .x(n90), .a(A[0]), .b(B[0]) );
	buf_2 U276 ( .x(n86), .a(A[31]) );
	buf_16 U277 ( .x(n88), .a(A[31]) );
	buf_16 U278 ( .x(n87), .a(A[31]) );
	nor2i_5 U279 ( .x(n126), .a(n127), .b(n128) );
	ao21_1 U28 ( .x(n296), .a(n170), .b(n247), .c(n128) );
	nor2_5 U280 ( .x(n165), .a(A[12]), .b(B[12]) );
	nor2i_3 U281 ( .x(n166), .a(n167), .b(n168) );
	exor2_3 U282 ( .x(SUM[5]), .a(n191), .b(n177) );
	exor2_3 U283 ( .x(SUM[29]), .a(n196), .b(n197) );
	exor2_3 U284 ( .x(SUM[26]), .a(n200), .b(n126) );
	exnor2_5 U285 ( .x(SUM[24]), .a(n166), .b(n203) );
	exnor2_3 U286 ( .x(SUM[23]), .a(n204), .b(n205) );
	exnor2_3 U287 ( .x(SUM[13]), .a(n107), .b(n144) );
	inv_6 U288 ( .x(n224), .a(B[15]) );
	nand2i_4 U289 ( .x(n225), .a(n165), .b(n226) );
	nand2i_3 U29 ( .x(n303), .a(n296), .b(n200) );
	oai211_4 U290 ( .x(n244), .a(n170), .b(n238), .c(n133), .d(n245) );
	oai21_5 U291 ( .x(n269), .a(n134), .b(n270), .c(n133) );
	exnor2_3 U292 ( .x(n272), .a(n269), .b(n88) );
	nor2i_5 U293 ( .x(n274), .a(n170), .b(n261) );
	aoi22_3 U294 ( .x(n259), .a(B[20]), .b(n88), .c(n87), .d(n264) );
	aoi21_3 U295 ( .x(n290), .a(n88), .b(n291), .c(n292) );
	nand2i_4 U296 ( .x(n293), .a(n251), .b(n294) );
	nand2_2 U297 ( .x(n297), .a(n253), .b(n255) );
	nand2i_4 U298 ( .x(n198), .a(n297), .b(n303) );
	inv_5 U299 ( .x(n168), .a(n262) );
	nand2_1 U30 ( .x(n255), .a(B[26]), .b(n87) );
	ao21_4 U300 ( .x(n195), .a(n208), .b(n311), .c(n313) );
	nand2i_4 U301 ( .x(n315), .a(B[7]), .b(n158) );
	oai211_4 U302 ( .x(n317), .a(n175), .b(n105), .c(n318), .d(n102) );
	nand2i_4 U303 ( .x(n319), .a(B[8]), .b(n220) );
	inv_5 U304 ( .x(n326), .a(n146) );
	nand2_5 U305 ( .x(n200), .a(n329), .b(n254) );
	aoai211_4 U306 ( .x(n196), .a(n52), .b(n329), .c(n170), .d(n333) );
	nand2i_4 U307 ( .x(n335), .a(n128), .b(n200) );
	nand2i_4 U308 ( .x(n199), .a(n322), .b(n335) );
	oai21_4 U309 ( .x(n205), .a(B[23]), .b(n88), .c(n300) );
	inv_2 U31 ( .x(n251), .a(B[28]) );
	inv_5 U310 ( .x(n270), .a(n211) );
	nand2_5 U311 ( .x(n341), .a(n339), .b(n315) );
	inv_5 U312 ( .x(n294), .a(n249) );
	or3i_5 U313 ( .x(n287), .a(n344), .b(n140), .c(n284) );
	nand2i_4 U314 ( .x(n288), .a(n142), .b(n327) );
	or3i_4 U315 ( .x(n340), .a(n192), .b(n103), .c(n277) );
	mux2i_3 U316 ( .x(n91), .d0(n276), .sl(n347), .d1(n272) );
	exor2_5 U317 ( .x(n203), .a(B[24]), .b(n87) );
	exor2_5 U318 ( .x(n197), .a(B[29]), .b(n88) );
	exor2_5 U319 ( .x(n194), .a(B[30]), .b(n88) );
	nand2i_0 U32 ( .x(n295), .a(n251), .b(n294) );
	exor2_5 U320 ( .x(n193), .a(B[31]), .b(n88) );
	nand2_8 U321 ( .x(n146), .a(n71), .b(A[12]) );
	inv_16 U322 ( .x(n170), .a(n87) );
	nand2i_6 U323 ( .x(n262), .a(n170), .b(n306) );
	aoi21_6 U324 ( .x(n120), .a(n121), .b(n122), .c(n87) );
	nand2_8 U325 ( .x(n254), .a(B[25]), .b(n88) );
	nor2i_6 U326 ( .x(n161), .a(n88), .b(n52) );
	nand2i_4 U327 ( .x(n331), .a(n170), .b(n82) );
	nand2i_5 U328 ( .x(n314), .a(B[4]), .b(n219) );
	nand2i_5 U329 ( .x(n231), .a(B[9]), .b(n221) );
	nand2_0 U33 ( .x(n127), .a(n50), .b(n87) );
	nand2i_5 U330 ( .x(n285), .a(A[14]), .b(n237) );
	nor2i_6 U331 ( .x(n122), .a(B[22]), .b(n223) );
	nand2i_5 U332 ( .x(n250), .a(n87), .b(n252) );
	nand2i_4 U333 ( .x(n339), .a(n157), .b(n340) );
	nand2i_4 U334 ( .x(n284), .a(n60), .b(n285) );
	exor2_2 U335 ( .x(SUM[20]), .a(n206), .b(n207) );
	inv_10 U336 ( .x(n184), .a(n171) );
	nand2i_4 U337 ( .x(n345), .a(n170), .b(n119) );
	mux2i_2 U338 ( .x(n96), .d0(n273), .sl(B[22]), .d1(n274) );
	exnor2_3 U339 ( .x(n273), .a(n261), .b(n170) );
	inv_1 U34 ( .x(n182), .a(n317) );
	nand2i_4 U340 ( .x(n59), .a(n72), .b(A[0]) );
	inv_0 U341 ( .x(n347), .a(n239) );
	inv_4 U342 ( .x(n68), .a(B[1]) );
	and2_4 U343 ( .x(n49), .a(A[1]), .b(B[1]) );
	inv_2 U35 ( .x(n215), .a(B[7]) );
	nand2i_2 U36 ( .x(n181), .a(n215), .b(n66) );
	nand2i_2 U37 ( .x(n180), .a(n158), .b(n66) );
	aoi21_1 U38 ( .x(n179), .a(n180), .b(n181), .c(n182) );
	inv_2 U39 ( .x(n234), .a(n71) );
	nand2i_2 U40 ( .x(n325), .a(A[12]), .b(n234) );
	inv_2 U41 ( .x(n238), .a(B[16]) );
	or3i_2 U42 ( .x(n241), .a(n242), .b(n238), .c(n239) );
	inv_2 U43 ( .x(n268), .a(n241) );
	ao21_1 U44 ( .x(n267), .a(n268), .b(n63), .c(n244) );
	inv_0 U45 ( .x(n118), .a(n264) );
	nand2i_3 U46 ( .x(n264), .a(n244), .b(n240) );
	nor2i_1 U47 ( .x(n132), .a(n133), .b(n134) );
	nand2_2 U48 ( .x(n133), .a(B[17]), .b(n86) );
	nand2i_2 U49 ( .x(n242), .a(n88), .b(n243) );
	exor2_2 U5 ( .x(SUM[30]), .a(n174), .b(n194) );
	inv_2 U50 ( .x(n243), .a(B[17]) );
	inv_2 U51 ( .x(n324), .a(n136) );
	nor2i_1 U52 ( .x(n148), .a(n85), .b(n150) );
	nand2i_2 U53 ( .x(n226), .a(B[11]), .b(n235) );
	nand2i_3 U54 ( .x(n261), .a(n183), .b(n262) );
	nor2_1 U56 ( .x(n298), .a(n260), .b(n223) );
	nand2_2 U57 ( .x(n299), .a(n263), .b(n300) );
	nand2i_4 U58 ( .x(n233), .a(n143), .b(n112) );
	inv_2 U59 ( .x(n112), .a(n227) );
	exnor2_3 U6 ( .x(SUM[31]), .a(n172), .b(n193) );
	or3i_4 U60 ( .x(n344), .a(n302), .b(n326), .c(n162) );
	nor2i_0 U61 ( .x(n101), .a(n102), .b(n103) );
	inv_2 U62 ( .x(n102), .a(n55) );
	and2_1 U63 ( .x(n55), .a(A[6]), .b(B[6]) );
	inv_5 U64 ( .x(n103), .a(n308) );
	aoai211_1 U65 ( .x(n190), .a(n217), .b(n218), .c(n321), .d(n178) );
	inv_2 U66 ( .x(n217), .a(A[5]) );
	inv_5 U67 ( .x(n218), .a(B[5]) );
	nand2_2 U68 ( .x(n142), .a(B[14]), .b(A[14]) );
	inv_5 U69 ( .x(n237), .a(B[14]) );
	aoi21_1 U70 ( .x(n111), .a(n112), .b(n109), .c(n113) );
	nand2i_2 U71 ( .x(n227), .a(n164), .b(n108) );
	nor2i_1 U72 ( .x(n113), .a(n159), .b(n160) );
	inv_0 U73 ( .x(n160), .a(n344) );
	inv_0 U74 ( .x(n153), .a(n280) );
	inv_2 U75 ( .x(n221), .a(A[9]) );
	nand2i_2 U76 ( .x(n229), .a(n230), .b(n231) );
	ao21_3 U77 ( .x(n208), .a(n312), .b(n70), .c(n49) );
	inv_2 U78 ( .x(n214), .a(B[2]) );
	inv_2 U79 ( .x(n252), .a(B[25]) );
	inv_0 U8 ( .x(n155), .a(n49) );
	nand2i_4 U80 ( .x(n291), .a(B[24]), .b(n278) );
	nor2i_5 U81 ( .x(n121), .a(B[24]), .b(n246) );
	inv_2 U82 ( .x(n246), .a(B[21]) );
	nor2i_0 U83 ( .x(n169), .a(n170), .b(n83) );
	exnor2_1 U84 ( .x(n275), .a(n83), .b(n170) );
	inv_2 U85 ( .x(n81), .a(n281) );
	inv_2 U86 ( .x(n286), .a(n288) );
	nand2i_2 U87 ( .x(n266), .a(n286), .b(n287) );
	nand2_2 U88 ( .x(n139), .a(B[15]), .b(n87) );
	inv_2 U89 ( .x(n134), .a(n242) );
	inv_2 U9 ( .x(n50), .a(n248) );
	nor2i_3 U90 ( .x(n276), .a(n269), .b(n87) );
	inv_2 U91 ( .x(n292), .a(n300) );
	nand2_2 U92 ( .x(n300), .a(B[23]), .b(n88) );
	inv_2 U93 ( .x(n223), .a(B[23]) );
	nand2_2 U94 ( .x(n263), .a(B[22]), .b(n88) );
	inv_2 U95 ( .x(n309), .a(n260) );
	nand2_2 U96 ( .x(n260), .a(B[21]), .b(B[22]) );
	nand2_2 U97 ( .x(n332), .a(B[29]), .b(n87) );
	inv_2 U98 ( .x(n222), .a(B[29]) );
	and4_4 U99 ( .x(n52), .a(n253), .b(n254), .c(n255), .d(n251) );

endmodule


module ID_test_1_desync (  INT, CLI, PIPEEMPTY, FREEZE, branch_address,
	branch_sig, Imm, rt_addr, rd_addr, reg_dst, reg_write, mem_to_reg, mem_write,
	mem_read, IR_opcode_field, IR_function_field, stall, counter, reset, NPC,
	IR_latched_input, reg_out_A, reg_out_B, reg_write_WB, WB_data, WB_data_old,
	test_si, test_so, test_se, sync_sel, global_g1, global_g2, Ctrl__Regs_1__en1,
	Ctrl__Regs_1__en2 );

input  INT, FREEZE, reset, reg_write_WB, test_si, test_se, sync_sel, global_g1,
	global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
input [31:0] NPC, IR_latched_input, WB_data, WB_data_old;
output  CLI, PIPEEMPTY, branch_sig, reg_dst, reg_write, mem_to_reg, mem_write,
	mem_read, stall, test_so;
output [1:0] counter;
output [31:0] branch_address, Imm, reg_out_A, reg_out_B;
output [4:0] rt_addr, rd_addr;
output [5:0] IR_opcode_field, IR_function_field;

wire CLI_reg__m2s, Cause_Reg_0, Cause_Reg_1, Cause_Reg_10, Cause_Reg_11,
	Cause_Reg_12, Cause_Reg_13, Cause_Reg_14, Cause_Reg_15, Cause_Reg_16,
	Cause_Reg_17, Cause_Reg_18, Cause_Reg_19, Cause_Reg_2, Cause_Reg_20, Cause_Reg_21,
	Cause_Reg_22, Cause_Reg_23, Cause_Reg_24, Cause_Reg_25, Cause_Reg_26,
	Cause_Reg_27, Cause_Reg_28, Cause_Reg_29, Cause_Reg_3, Cause_Reg_30, Cause_Reg_31,
	Cause_Reg_4, Cause_Reg_5, Cause_Reg_6, Cause_Reg_7, Cause_Reg_8, Cause_Reg_9,
	Cause_Reg_reg_0__m2s, Cause_Reg_reg_10__m2s, Cause_Reg_reg_11__m2s, Cause_Reg_reg_12__m2s,
	Cause_Reg_reg_13__m2s, Cause_Reg_reg_14__m2s, Cause_Reg_reg_15__m2s, Cause_Reg_reg_16__m2s,
	Cause_Reg_reg_17__m2s, Cause_Reg_reg_18__m2s, Cause_Reg_reg_19__m2s, Cause_Reg_reg_1__m2s,
	Cause_Reg_reg_20__m2s, Cause_Reg_reg_21__m2s, Cause_Reg_reg_22__m2s, Cause_Reg_reg_23__m2s,
	Cause_Reg_reg_24__m2s, Cause_Reg_reg_25__m2s, Cause_Reg_reg_26__m2s, Cause_Reg_reg_27__m2s,
	Cause_Reg_reg_28__m2s, Cause_Reg_reg_29__m2s, Cause_Reg_reg_2__m2s, Cause_Reg_reg_30__m2s,
	Cause_Reg_reg_31__m2s, Cause_Reg_reg_3__m2s, Cause_Reg_reg_4__m2s, Cause_Reg_reg_5__m2s,
	Cause_Reg_reg_6__m2s, Cause_Reg_reg_7__m2s, Cause_Reg_reg_8__m2s, Cause_Reg_reg_9__m2s,
	EPC_0, EPC_1, EPC_10, EPC_11, EPC_12, EPC_13, EPC_14, EPC_15, EPC_16,
	EPC_17, EPC_18, EPC_19, EPC_2, EPC_20, EPC_21, EPC_22, EPC_23, EPC_24,
	EPC_25, EPC_26, EPC_27, EPC_28, EPC_29, EPC_3, EPC_30, EPC_31, EPC_4,
	EPC_5, EPC_6, EPC_7, EPC_8, EPC_9, EPC_reg_0__m2s, EPC_reg_10__m2s, EPC_reg_11__m2s,
	EPC_reg_12__m2s, EPC_reg_13__m2s, EPC_reg_14__m2s, EPC_reg_15__m2s, EPC_reg_16__m2s,
	EPC_reg_17__m2s, EPC_reg_18__m2s, EPC_reg_19__m2s, EPC_reg_1__m2s, EPC_reg_20__m2s,
	EPC_reg_21__m2s, EPC_reg_22__m2s, EPC_reg_23__m2s, EPC_reg_24__m2s, EPC_reg_25__m2s,
	EPC_reg_26__m2s, EPC_reg_27__m2s, EPC_reg_28__m2s, EPC_reg_29__m2s, EPC_reg_2__m2s,
	EPC_reg_30__m2s, EPC_reg_31__m2s, EPC_reg_3__m2s, EPC_reg_4__m2s, EPC_reg_5__m2s,
	EPC_reg_6__m2s, EPC_reg_7__m2s, EPC_reg_8__m2s, EPC_reg_9__m2s, IR_function_field_reg_0__m2s,
	IR_function_field_reg_1__m2s, IR_function_field_reg_2__m2s, IR_function_field_reg_3__m2s,
	IR_function_field_reg_4__m2s, IR_function_field_reg_5__m2s, IR_latched_0,
	IR_latched_1, IR_latched_10, IR_latched_11, IR_latched_12, IR_latched_13,
	IR_latched_14, IR_latched_15, IR_latched_2, IR_latched_3, IR_latched_4,
	IR_latched_5, IR_latched_8, IR_latched_9, IR_opcode_field_reg_0__m2s,
	IR_opcode_field_reg_1__m2s, IR_opcode_field_reg_2__m2s, IR_opcode_field_reg_3__m2s,
	IR_opcode_field_reg_4__m2s, IR_opcode_field_reg_5__m2s, Imm_reg_0__m2s,
	Imm_reg_10__m2s, Imm_reg_11__m2s, Imm_reg_12__m2s, Imm_reg_13__m2s, Imm_reg_14__m2s,
	Imm_reg_15__m2s, Imm_reg_16__m2s, Imm_reg_17__m2s, Imm_reg_18__m2s, Imm_reg_19__m2s,
	Imm_reg_1__m2s, Imm_reg_20__m2s, Imm_reg_21__m2s, Imm_reg_22__m2s, Imm_reg_23__m2s,
	Imm_reg_24__m2s, Imm_reg_25__m2s, Imm_reg_26__m2s, Imm_reg_27__m2s, Imm_reg_28__m2s,
	Imm_reg_29__m2s, Imm_reg_2__m2s, Imm_reg_30__m2s, Imm_reg_31__m2s, Imm_reg_3__m2s,
	Imm_reg_4__m2s, Imm_reg_5__m2s, Imm_reg_6__m2s, Imm_reg_7__m2s, Imm_reg_8__m2s,
	Imm_reg_9__m2s, N13832, N437, N438, N439, N440, N441, N442, N443, N444,
	N445, N446, N447, N448, N449, N450, N451, N452, N453, N454, N455, N456,
	N457, N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
	N504, N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
	N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526, N527,
	N528, N529, N530, N531, N5319, N532, N5320, N5321, N5322, N5323, N5324,
	N5325, N5326, N5327, N5328, N5329, N533, N5330, N5331, N5332, N5333, N5334,
	N5335, N5336, N5337, N5338, N5339, N534, N5340, N5341, N5342, N5343, N5344,
	N5345, N5346, N5347, N5348, N5349, N535, N5350, N5351, N5352, N5353, N5354,
	N5355, N5356, N5357, N5358, N5359, N5360, N5361, N5362, N5363, N5364,
	N5365, N5366, N5367, N5368, N5369, N5370, N5371, N5372, N5373, N5374,
	N5375, N5376, N5377, N5378, N5379, N5380, N5381, N5382, N5387, N5388,
	N5389, N5390, N5391, N5392, N5393, N5394, N5395, N5396, N5397, N5398,
	N5399, N5400, N5401, N5402, N5403, N5404, N5405, N5406, N5407, N5408,
	N5409, N5410, N5411, N5412, N5413, N5414, N5415, N5416, N5417, N5418,
	N5419, N5420, N5421, N5422, N5423, N5424, N5425, N5426, N5427, N5428,
	N5429, N5430, N5431, N5432, N5433, N5434, N5435, N5436, N5437, N5438,
	N5439, N5440, N5441, N5442, N5443, N5444, N5445, N5446, N5447, N5448,
	N5449, N5450, N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993,
	N5994, N5995, N5996, N5997, N5998, N5999, N6000, N6001, N6002, N6003,
	N6004, N6005, N6006, N6007, N6008, N6009, N6010, N6011, N6012, N6013,
	N6014, N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022, N6023,
	N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032, N6033,
	N6034, N6035, N6036, N6037, N6038, N6039, N6040, N6041, N6042, N6043,
	N6044, N6045, N6046, N6047, N6048, N6049, N6328, N6332, N6334, N6336,
	N6338, N6340, N6342, N6344, N6346, N6348, N6350, N6352, N6354, N6356,
	N6358, N6360, N6362, N6364, N6366, N6368, N6370, N6376, N6380, N6382,
	N6384, N6386, N6388, N6390, N6718, N6719, N6720, N6721, N6722, N6723,
	N6724, N6725, N6726, N6727, N6728, N6729, N6730, N6731, N6732, N6733,
	N6734, N6735, N6736, N6737, N6738, N6739, N6740, N6741, N6742, N6743,
	N6744, N6745, N6746, N6747, N6748, N6749, WB_index_0, WB_index_1, WB_index_2,
	WB_index_3, WB_index_4, WB_index_reg_0__m2s, WB_index_reg_1__m2s, WB_index_reg_2__m2s,
	WB_index_reg_3__m2s, WB_index_reg_4__m2s, _EPC_reg_31_net69891, _RegFile_0__0,
	_RegFile_0__1, _RegFile_0__10, _RegFile_0__11, _RegFile_0__12, _RegFile_0__13,
	_RegFile_0__14, _RegFile_0__15, _RegFile_0__16, _RegFile_0__17, _RegFile_0__18,
	_RegFile_0__19, _RegFile_0__2, _RegFile_0__20, _RegFile_0__21, _RegFile_0__22,
	_RegFile_0__23, _RegFile_0__24, _RegFile_0__25, _RegFile_0__26, _RegFile_0__27,
	_RegFile_0__28, _RegFile_0__29, _RegFile_0__3, _RegFile_0__30, _RegFile_0__31,
	_RegFile_0__4, _RegFile_0__5, _RegFile_0__6, _RegFile_0__7, _RegFile_0__8,
	_RegFile_0__9, _RegFile_10__0, _RegFile_10__1, _RegFile_10__10, _RegFile_10__11,
	_RegFile_10__12, _RegFile_10__13, _RegFile_10__14, _RegFile_10__15, _RegFile_10__16,
	_RegFile_10__17, _RegFile_10__18, _RegFile_10__19, _RegFile_10__2, _RegFile_10__20,
	_RegFile_10__21, _RegFile_10__22, _RegFile_10__23, _RegFile_10__24, _RegFile_10__25,
	_RegFile_10__26, _RegFile_10__27, _RegFile_10__28, _RegFile_10__29, _RegFile_10__3,
	_RegFile_10__30, _RegFile_10__31, _RegFile_10__4, _RegFile_10__5, _RegFile_10__6,
	_RegFile_10__7, _RegFile_10__8, _RegFile_10__9, _RegFile_11__0, _RegFile_11__1,
	_RegFile_11__10, _RegFile_11__11, _RegFile_11__12, _RegFile_11__13, _RegFile_11__14,
	_RegFile_11__15, _RegFile_11__16, _RegFile_11__17, _RegFile_11__18, _RegFile_11__19,
	_RegFile_11__2, _RegFile_11__20, _RegFile_11__21, _RegFile_11__22, _RegFile_11__23,
	_RegFile_11__24, _RegFile_11__25, _RegFile_11__26, _RegFile_11__27, _RegFile_11__28,
	_RegFile_11__29, _RegFile_11__3, _RegFile_11__30, _RegFile_11__31, _RegFile_11__4,
	_RegFile_11__5, _RegFile_11__6, _RegFile_11__7, _RegFile_11__8, _RegFile_11__9,
	_RegFile_12__0, _RegFile_12__1, _RegFile_12__10, _RegFile_12__11, _RegFile_12__12,
	_RegFile_12__13, _RegFile_12__14, _RegFile_12__15, _RegFile_12__16, _RegFile_12__17,
	_RegFile_12__18, _RegFile_12__19, _RegFile_12__2, _RegFile_12__20, _RegFile_12__21,
	_RegFile_12__22, _RegFile_12__23, _RegFile_12__24, _RegFile_12__25, _RegFile_12__26,
	_RegFile_12__27, _RegFile_12__28, _RegFile_12__29, _RegFile_12__3, _RegFile_12__30,
	_RegFile_12__31, _RegFile_12__4, _RegFile_12__5, _RegFile_12__6, _RegFile_12__7,
	_RegFile_12__8, _RegFile_12__9, _RegFile_13__0, _RegFile_13__1, _RegFile_13__10,
	_RegFile_13__11, _RegFile_13__12, _RegFile_13__13, _RegFile_13__14, _RegFile_13__15,
	_RegFile_13__16, _RegFile_13__17, _RegFile_13__18, _RegFile_13__19, _RegFile_13__2,
	_RegFile_13__20, _RegFile_13__21, _RegFile_13__22, _RegFile_13__23, _RegFile_13__24,
	_RegFile_13__25, _RegFile_13__26, _RegFile_13__27, _RegFile_13__28, _RegFile_13__29,
	_RegFile_13__3, _RegFile_13__30, _RegFile_13__31, _RegFile_13__4, _RegFile_13__5,
	_RegFile_13__6, _RegFile_13__7, _RegFile_13__8, _RegFile_13__9, _RegFile_14__0,
	_RegFile_14__1, _RegFile_14__10, _RegFile_14__11, _RegFile_14__12, _RegFile_14__13,
	_RegFile_14__14, _RegFile_14__15, _RegFile_14__16, _RegFile_14__17, _RegFile_14__18,
	_RegFile_14__19, _RegFile_14__2, _RegFile_14__20, _RegFile_14__21, _RegFile_14__22,
	_RegFile_14__23, _RegFile_14__24, _RegFile_14__25, _RegFile_14__26, _RegFile_14__27,
	_RegFile_14__28, _RegFile_14__29, _RegFile_14__3, _RegFile_14__30, _RegFile_14__31,
	_RegFile_14__4, _RegFile_14__5, _RegFile_14__6, _RegFile_14__7, _RegFile_14__8,
	_RegFile_14__9, _RegFile_15__0, _RegFile_15__1, _RegFile_15__10, _RegFile_15__11,
	_RegFile_15__12, _RegFile_15__13, _RegFile_15__14, _RegFile_15__15, _RegFile_15__16,
	_RegFile_15__17, _RegFile_15__18, _RegFile_15__19, _RegFile_15__2, _RegFile_15__20,
	_RegFile_15__21, _RegFile_15__22, _RegFile_15__23, _RegFile_15__24, _RegFile_15__25,
	_RegFile_15__26, _RegFile_15__27, _RegFile_15__28, _RegFile_15__29, _RegFile_15__3,
	_RegFile_15__30, _RegFile_15__31, _RegFile_15__4, _RegFile_15__5, _RegFile_15__6,
	_RegFile_15__7, _RegFile_15__8, _RegFile_15__9, _RegFile_16__0, _RegFile_16__1,
	_RegFile_16__10, _RegFile_16__11, _RegFile_16__12, _RegFile_16__13, _RegFile_16__14,
	_RegFile_16__15, _RegFile_16__16, _RegFile_16__17, _RegFile_16__18, _RegFile_16__19,
	_RegFile_16__2, _RegFile_16__20, _RegFile_16__21, _RegFile_16__22, _RegFile_16__23,
	_RegFile_16__24, _RegFile_16__25, _RegFile_16__26, _RegFile_16__27, _RegFile_16__28,
	_RegFile_16__29, _RegFile_16__3, _RegFile_16__30, _RegFile_16__31, _RegFile_16__4,
	_RegFile_16__5, _RegFile_16__6, _RegFile_16__7, _RegFile_16__8, _RegFile_16__9,
	_RegFile_17__0, _RegFile_17__1, _RegFile_17__10, _RegFile_17__11, _RegFile_17__12,
	_RegFile_17__13, _RegFile_17__14, _RegFile_17__15, _RegFile_17__16, _RegFile_17__17,
	_RegFile_17__18, _RegFile_17__19, _RegFile_17__2, _RegFile_17__20, _RegFile_17__21,
	_RegFile_17__22, _RegFile_17__23, _RegFile_17__24, _RegFile_17__25, _RegFile_17__26,
	_RegFile_17__27, _RegFile_17__28, _RegFile_17__29, _RegFile_17__3, _RegFile_17__30,
	_RegFile_17__31, _RegFile_17__4, _RegFile_17__5, _RegFile_17__6, _RegFile_17__7,
	_RegFile_17__8, _RegFile_17__9, _RegFile_18__0, _RegFile_18__1, _RegFile_18__10,
	_RegFile_18__11, _RegFile_18__12, _RegFile_18__13, _RegFile_18__14, _RegFile_18__15,
	_RegFile_18__16, _RegFile_18__17, _RegFile_18__18, _RegFile_18__19, _RegFile_18__2,
	_RegFile_18__20, _RegFile_18__21, _RegFile_18__22, _RegFile_18__23, _RegFile_18__24,
	_RegFile_18__25, _RegFile_18__26, _RegFile_18__27, _RegFile_18__28, _RegFile_18__29,
	_RegFile_18__3, _RegFile_18__30, _RegFile_18__31, _RegFile_18__4, _RegFile_18__5,
	_RegFile_18__6, _RegFile_18__7, _RegFile_18__8, _RegFile_18__9, _RegFile_19__0,
	_RegFile_19__1, _RegFile_19__10, _RegFile_19__11, _RegFile_19__12, _RegFile_19__13,
	_RegFile_19__14, _RegFile_19__15, _RegFile_19__16, _RegFile_19__17, _RegFile_19__18,
	_RegFile_19__19, _RegFile_19__2, _RegFile_19__20, _RegFile_19__21, _RegFile_19__22,
	_RegFile_19__23, _RegFile_19__24, _RegFile_19__25, _RegFile_19__26, _RegFile_19__27,
	_RegFile_19__28, _RegFile_19__29, _RegFile_19__3, _RegFile_19__30, _RegFile_19__31,
	_RegFile_19__4, _RegFile_19__5, _RegFile_19__6, _RegFile_19__7, _RegFile_19__8,
	_RegFile_19__9, _RegFile_1__0, _RegFile_1__1, _RegFile_1__10, _RegFile_1__11,
	_RegFile_1__12, _RegFile_1__13, _RegFile_1__14, _RegFile_1__15, _RegFile_1__16,
	_RegFile_1__17, _RegFile_1__18, _RegFile_1__19, _RegFile_1__2, _RegFile_1__20,
	_RegFile_1__21, _RegFile_1__22, _RegFile_1__23, _RegFile_1__24, _RegFile_1__25,
	_RegFile_1__26, _RegFile_1__27, _RegFile_1__28, _RegFile_1__29, _RegFile_1__3,
	_RegFile_1__30, _RegFile_1__31, _RegFile_1__4, _RegFile_1__5, _RegFile_1__6,
	_RegFile_1__7, _RegFile_1__8, _RegFile_1__9, _RegFile_20__0, _RegFile_20__1,
	_RegFile_20__10, _RegFile_20__11, _RegFile_20__12, _RegFile_20__13, _RegFile_20__14,
	_RegFile_20__15, _RegFile_20__16, _RegFile_20__17, _RegFile_20__18, _RegFile_20__19,
	_RegFile_20__2, _RegFile_20__20, _RegFile_20__21, _RegFile_20__22, _RegFile_20__23,
	_RegFile_20__24, _RegFile_20__25, _RegFile_20__26, _RegFile_20__27, _RegFile_20__28,
	_RegFile_20__29, _RegFile_20__3, _RegFile_20__30, _RegFile_20__31, _RegFile_20__4,
	_RegFile_20__5, _RegFile_20__6, _RegFile_20__7, _RegFile_20__8, _RegFile_20__9,
	_RegFile_21__0, _RegFile_21__1, _RegFile_21__10, _RegFile_21__11, _RegFile_21__12,
	_RegFile_21__13, _RegFile_21__14, _RegFile_21__15, _RegFile_21__16, _RegFile_21__17,
	_RegFile_21__18, _RegFile_21__19, _RegFile_21__2, _RegFile_21__20, _RegFile_21__21,
	_RegFile_21__22, _RegFile_21__23, _RegFile_21__24, _RegFile_21__25, _RegFile_21__26,
	_RegFile_21__27, _RegFile_21__28, _RegFile_21__29, _RegFile_21__3, _RegFile_21__30,
	_RegFile_21__31, _RegFile_21__4, _RegFile_21__5, _RegFile_21__6, _RegFile_21__7,
	_RegFile_21__8, _RegFile_21__9, _RegFile_22__0, _RegFile_22__1, _RegFile_22__10,
	_RegFile_22__11, _RegFile_22__12, _RegFile_22__13, _RegFile_22__14, _RegFile_22__15,
	_RegFile_22__16, _RegFile_22__17, _RegFile_22__18, _RegFile_22__19, _RegFile_22__2,
	_RegFile_22__20, _RegFile_22__21, _RegFile_22__22, _RegFile_22__23, _RegFile_22__24,
	_RegFile_22__25, _RegFile_22__26, _RegFile_22__27, _RegFile_22__28, _RegFile_22__29,
	_RegFile_22__3, _RegFile_22__30, _RegFile_22__31, _RegFile_22__4, _RegFile_22__5,
	_RegFile_22__6, _RegFile_22__7, _RegFile_22__8, _RegFile_22__9, _RegFile_23__0,
	_RegFile_23__1, _RegFile_23__10, _RegFile_23__11, _RegFile_23__12, _RegFile_23__13,
	_RegFile_23__14, _RegFile_23__15, _RegFile_23__16, _RegFile_23__17, _RegFile_23__18,
	_RegFile_23__19, _RegFile_23__2, _RegFile_23__20, _RegFile_23__21, _RegFile_23__22,
	_RegFile_23__23, _RegFile_23__24, _RegFile_23__25, _RegFile_23__26, _RegFile_23__27,
	_RegFile_23__28, _RegFile_23__29, _RegFile_23__3, _RegFile_23__30, _RegFile_23__31,
	_RegFile_23__4, _RegFile_23__5, _RegFile_23__6, _RegFile_23__7, _RegFile_23__8,
	_RegFile_23__9, _RegFile_24__0, _RegFile_24__1, _RegFile_24__10, _RegFile_24__11,
	_RegFile_24__12, _RegFile_24__13, _RegFile_24__14, _RegFile_24__15, _RegFile_24__16,
	_RegFile_24__17, _RegFile_24__18, _RegFile_24__19, _RegFile_24__2, _RegFile_24__20,
	_RegFile_24__21, _RegFile_24__22, _RegFile_24__23, _RegFile_24__24, _RegFile_24__25,
	_RegFile_24__26, _RegFile_24__27, _RegFile_24__28, _RegFile_24__29, _RegFile_24__3,
	_RegFile_24__30, _RegFile_24__31, _RegFile_24__4, _RegFile_24__5, _RegFile_24__6,
	_RegFile_24__7, _RegFile_24__8, _RegFile_24__9, _RegFile_25__0, _RegFile_25__1,
	_RegFile_25__10, _RegFile_25__11, _RegFile_25__12, _RegFile_25__13, _RegFile_25__14,
	_RegFile_25__15, _RegFile_25__16, _RegFile_25__17, _RegFile_25__18, _RegFile_25__19,
	_RegFile_25__2, _RegFile_25__20, _RegFile_25__21, _RegFile_25__22, _RegFile_25__23,
	_RegFile_25__24, _RegFile_25__25, _RegFile_25__26, _RegFile_25__27, _RegFile_25__28,
	_RegFile_25__29, _RegFile_25__3, _RegFile_25__30, _RegFile_25__31, _RegFile_25__4,
	_RegFile_25__5, _RegFile_25__6, _RegFile_25__7, _RegFile_25__8, _RegFile_25__9,
	_RegFile_26__0, _RegFile_26__1, _RegFile_26__10, _RegFile_26__11, _RegFile_26__12,
	_RegFile_26__13, _RegFile_26__14, _RegFile_26__15, _RegFile_26__16, _RegFile_26__17,
	_RegFile_26__18, _RegFile_26__19, _RegFile_26__2, _RegFile_26__20, _RegFile_26__21,
	_RegFile_26__22, _RegFile_26__23, _RegFile_26__24, _RegFile_26__25, _RegFile_26__26,
	_RegFile_26__27, _RegFile_26__28, _RegFile_26__29, _RegFile_26__3, _RegFile_26__30,
	_RegFile_26__31, _RegFile_26__4, _RegFile_26__5, _RegFile_26__6, _RegFile_26__7,
	_RegFile_26__8, _RegFile_26__9, _RegFile_27__0, _RegFile_27__1, _RegFile_27__10,
	_RegFile_27__11, _RegFile_27__12, _RegFile_27__13, _RegFile_27__14, _RegFile_27__15,
	_RegFile_27__16, _RegFile_27__17, _RegFile_27__18, _RegFile_27__19, _RegFile_27__2,
	_RegFile_27__20, _RegFile_27__21, _RegFile_27__22, _RegFile_27__23, _RegFile_27__24,
	_RegFile_27__25, _RegFile_27__26, _RegFile_27__27, _RegFile_27__28, _RegFile_27__29,
	_RegFile_27__3, _RegFile_27__30, _RegFile_27__31, _RegFile_27__4, _RegFile_27__5,
	_RegFile_27__6, _RegFile_27__7, _RegFile_27__8, _RegFile_27__9, _RegFile_28__0,
	_RegFile_28__1, _RegFile_28__10, _RegFile_28__11, _RegFile_28__12, _RegFile_28__13,
	_RegFile_28__14, _RegFile_28__15, _RegFile_28__16, _RegFile_28__17, _RegFile_28__18,
	_RegFile_28__19, _RegFile_28__2, _RegFile_28__20, _RegFile_28__21, _RegFile_28__22,
	_RegFile_28__23, _RegFile_28__24, _RegFile_28__25, _RegFile_28__26, _RegFile_28__27,
	_RegFile_28__28, _RegFile_28__29, _RegFile_28__3, _RegFile_28__30, _RegFile_28__31,
	_RegFile_28__4, _RegFile_28__5, _RegFile_28__6, _RegFile_28__7, _RegFile_28__8,
	_RegFile_28__9, _RegFile_29__0, _RegFile_29__1, _RegFile_29__10, _RegFile_29__11,
	_RegFile_29__12, _RegFile_29__13, _RegFile_29__14, _RegFile_29__15, _RegFile_29__16,
	_RegFile_29__17, _RegFile_29__18, _RegFile_29__19, _RegFile_29__2, _RegFile_29__20,
	_RegFile_29__21, _RegFile_29__22, _RegFile_29__23, _RegFile_29__24, _RegFile_29__25,
	_RegFile_29__26, _RegFile_29__27, _RegFile_29__28, _RegFile_29__29, _RegFile_29__3,
	_RegFile_29__30, _RegFile_29__31, _RegFile_29__4, _RegFile_29__5, _RegFile_29__6,
	_RegFile_29__7, _RegFile_29__8, _RegFile_29__9, _RegFile_2__0, _RegFile_2__1,
	_RegFile_2__10, _RegFile_2__11, _RegFile_2__12, _RegFile_2__13, _RegFile_2__14,
	_RegFile_2__15, _RegFile_2__16, _RegFile_2__17, _RegFile_2__18, _RegFile_2__19,
	_RegFile_2__2, _RegFile_2__20, _RegFile_2__21, _RegFile_2__22, _RegFile_2__23,
	_RegFile_2__24, _RegFile_2__25, _RegFile_2__26, _RegFile_2__27, _RegFile_2__28,
	_RegFile_2__29, _RegFile_2__3, _RegFile_2__30, _RegFile_2__31, _RegFile_2__4,
	_RegFile_2__5, _RegFile_2__6, _RegFile_2__7, _RegFile_2__8, _RegFile_2__9,
	_RegFile_30__0, _RegFile_30__1, _RegFile_30__10, _RegFile_30__11, _RegFile_30__12,
	_RegFile_30__13, _RegFile_30__14, _RegFile_30__15, _RegFile_30__16, _RegFile_30__17,
	_RegFile_30__18, _RegFile_30__19, _RegFile_30__2, _RegFile_30__20, _RegFile_30__21,
	_RegFile_30__22, _RegFile_30__23, _RegFile_30__24, _RegFile_30__25, _RegFile_30__26,
	_RegFile_30__27, _RegFile_30__28, _RegFile_30__29, _RegFile_30__3, _RegFile_30__30,
	_RegFile_30__31, _RegFile_30__4, _RegFile_30__5, _RegFile_30__6, _RegFile_30__7,
	_RegFile_30__8, _RegFile_30__9, _RegFile_31__0, _RegFile_31__1, _RegFile_31__10,
	_RegFile_31__11, _RegFile_31__12, _RegFile_31__13, _RegFile_31__14, _RegFile_31__15,
	_RegFile_31__16, _RegFile_31__17, _RegFile_31__18, _RegFile_31__19, _RegFile_31__2,
	_RegFile_31__20, _RegFile_31__21, _RegFile_31__22, _RegFile_31__23, _RegFile_31__24,
	_RegFile_31__25, _RegFile_31__26, _RegFile_31__27, _RegFile_31__28, _RegFile_31__29,
	_RegFile_31__3, _RegFile_31__30, _RegFile_31__31, _RegFile_31__4, _RegFile_31__5,
	_RegFile_31__6, _RegFile_31__7, _RegFile_31__8, _RegFile_31__9, _RegFile_3__0,
	_RegFile_3__1, _RegFile_3__10, _RegFile_3__11, _RegFile_3__12, _RegFile_3__13,
	_RegFile_3__14, _RegFile_3__15, _RegFile_3__16, _RegFile_3__17, _RegFile_3__18,
	_RegFile_3__19, _RegFile_3__2, _RegFile_3__20, _RegFile_3__21, _RegFile_3__22,
	_RegFile_3__23, _RegFile_3__24, _RegFile_3__25, _RegFile_3__26, _RegFile_3__27,
	_RegFile_3__28, _RegFile_3__29, _RegFile_3__3, _RegFile_3__30, _RegFile_3__31,
	_RegFile_3__4, _RegFile_3__5, _RegFile_3__6, _RegFile_3__7, _RegFile_3__8,
	_RegFile_3__9, _RegFile_4__0, _RegFile_4__1, _RegFile_4__10, _RegFile_4__11,
	_RegFile_4__12, _RegFile_4__13, _RegFile_4__14, _RegFile_4__15, _RegFile_4__16,
	_RegFile_4__17, _RegFile_4__18, _RegFile_4__19, _RegFile_4__2, _RegFile_4__20,
	_RegFile_4__21, _RegFile_4__22, _RegFile_4__23, _RegFile_4__24, _RegFile_4__25,
	_RegFile_4__26, _RegFile_4__27, _RegFile_4__28, _RegFile_4__29, _RegFile_4__3,
	_RegFile_4__30, _RegFile_4__31, _RegFile_4__4, _RegFile_4__5, _RegFile_4__6,
	_RegFile_4__7, _RegFile_4__8, _RegFile_4__9, _RegFile_5__0, _RegFile_5__1,
	_RegFile_5__10, _RegFile_5__11, _RegFile_5__12, _RegFile_5__13, _RegFile_5__14,
	_RegFile_5__15, _RegFile_5__16, _RegFile_5__17, _RegFile_5__18, _RegFile_5__19,
	_RegFile_5__2, _RegFile_5__20, _RegFile_5__21, _RegFile_5__22, _RegFile_5__23,
	_RegFile_5__24, _RegFile_5__25, _RegFile_5__26, _RegFile_5__27, _RegFile_5__28,
	_RegFile_5__29, _RegFile_5__3, _RegFile_5__30, _RegFile_5__31, _RegFile_5__4,
	_RegFile_5__5, _RegFile_5__6, _RegFile_5__7, _RegFile_5__8, _RegFile_5__9,
	_RegFile_6__0, _RegFile_6__1, _RegFile_6__10, _RegFile_6__11, _RegFile_6__12,
	_RegFile_6__13, _RegFile_6__14, _RegFile_6__15, _RegFile_6__16, _RegFile_6__17,
	_RegFile_6__18, _RegFile_6__19, _RegFile_6__2, _RegFile_6__20, _RegFile_6__21,
	_RegFile_6__22, _RegFile_6__23, _RegFile_6__24, _RegFile_6__25, _RegFile_6__26,
	_RegFile_6__27, _RegFile_6__28, _RegFile_6__29, _RegFile_6__3, _RegFile_6__30,
	_RegFile_6__31, _RegFile_6__4, _RegFile_6__5, _RegFile_6__6, _RegFile_6__7,
	_RegFile_6__8, _RegFile_6__9, _RegFile_7__0, _RegFile_7__1, _RegFile_7__10,
	_RegFile_7__11, _RegFile_7__12, _RegFile_7__13, _RegFile_7__14, _RegFile_7__15,
	_RegFile_7__16, _RegFile_7__17, _RegFile_7__18, _RegFile_7__19, _RegFile_7__2,
	_RegFile_7__20, _RegFile_7__21, _RegFile_7__22, _RegFile_7__23, _RegFile_7__24,
	_RegFile_7__25, _RegFile_7__26, _RegFile_7__27, _RegFile_7__28, _RegFile_7__29,
	_RegFile_7__3, _RegFile_7__30, _RegFile_7__31, _RegFile_7__4, _RegFile_7__5,
	_RegFile_7__6, _RegFile_7__7, _RegFile_7__8, _RegFile_7__9, _RegFile_8__0,
	_RegFile_8__1, _RegFile_8__10, _RegFile_8__11, _RegFile_8__12, _RegFile_8__13,
	_RegFile_8__14, _RegFile_8__15, _RegFile_8__16, _RegFile_8__17, _RegFile_8__18,
	_RegFile_8__19, _RegFile_8__2, _RegFile_8__20, _RegFile_8__21, _RegFile_8__22,
	_RegFile_8__23, _RegFile_8__24, _RegFile_8__25, _RegFile_8__26, _RegFile_8__27,
	_RegFile_8__28, _RegFile_8__29, _RegFile_8__3, _RegFile_8__30, _RegFile_8__31,
	_RegFile_8__4, _RegFile_8__5, _RegFile_8__6, _RegFile_8__7, _RegFile_8__8,
	_RegFile_8__9, _RegFile_9__0, _RegFile_9__1, _RegFile_9__10, _RegFile_9__11,
	_RegFile_9__12, _RegFile_9__13, _RegFile_9__14, _RegFile_9__15, _RegFile_9__16,
	_RegFile_9__17, _RegFile_9__18, _RegFile_9__19, _RegFile_9__2, _RegFile_9__20,
	_RegFile_9__21, _RegFile_9__22, _RegFile_9__23, _RegFile_9__24, _RegFile_9__25,
	_RegFile_9__26, _RegFile_9__27, _RegFile_9__28, _RegFile_9__29, _RegFile_9__3,
	_RegFile_9__30, _RegFile_9__31, _RegFile_9__4, _RegFile_9__5, _RegFile_9__6,
	_RegFile_9__7, _RegFile_9__8, _RegFile_9__9, _RegFile_reg_0__0__m2s, _RegFile_reg_0__10__m2s,
	_RegFile_reg_0__11__m2s, _RegFile_reg_0__12__m2s, _RegFile_reg_0__13__m2s,
	_RegFile_reg_0__14__m2s, _RegFile_reg_0__15__m2s, _RegFile_reg_0__16__m2s,
	_RegFile_reg_0__17__m2s, _RegFile_reg_0__18__m2s, _RegFile_reg_0__19__m2s,
	_RegFile_reg_0__1__m2s, _RegFile_reg_0__20__m2s, _RegFile_reg_0__21__m2s,
	_RegFile_reg_0__22__m2s, _RegFile_reg_0__23__m2s, _RegFile_reg_0__24__m2s,
	_RegFile_reg_0__25__m2s, _RegFile_reg_0__26__m2s, _RegFile_reg_0__27__m2s,
	_RegFile_reg_0__28__m2s, _RegFile_reg_0__29__m2s, _RegFile_reg_0__2__m2s,
	_RegFile_reg_0__30__m2s, _RegFile_reg_0__31__m2s, _RegFile_reg_0__3__m2s,
	_RegFile_reg_0__4__m2s, _RegFile_reg_0__5__m2s, _RegFile_reg_0__6__m2s,
	_RegFile_reg_0__7__m2s, _RegFile_reg_0__8__m2s, _RegFile_reg_0__9__m2s,
	_RegFile_reg_10__0__m2s, _RegFile_reg_10__10__m2s, _RegFile_reg_10__11__m2s,
	_RegFile_reg_10__12__m2s, _RegFile_reg_10__13__m2s, _RegFile_reg_10__14__m2s,
	_RegFile_reg_10__15__m2s, _RegFile_reg_10__16__m2s, _RegFile_reg_10__17__m2s,
	_RegFile_reg_10__18__m2s, _RegFile_reg_10__19__m2s, _RegFile_reg_10__1__m2s,
	_RegFile_reg_10__20__m2s, _RegFile_reg_10__21__m2s, _RegFile_reg_10__22__m2s,
	_RegFile_reg_10__23__m2s, _RegFile_reg_10__24__m2s, _RegFile_reg_10__25__m2s,
	_RegFile_reg_10__26__m2s, _RegFile_reg_10__27__m2s, _RegFile_reg_10__28__m2s,
	_RegFile_reg_10__29__m2s, _RegFile_reg_10__2__m2s, _RegFile_reg_10__30__m2s,
	_RegFile_reg_10__31__m2s, _RegFile_reg_10__3__m2s, _RegFile_reg_10__4__m2s,
	_RegFile_reg_10__5__m2s, _RegFile_reg_10__6__m2s, _RegFile_reg_10__7__m2s,
	_RegFile_reg_10__8__m2s, _RegFile_reg_10__9__m2s, _RegFile_reg_11__0__m2s,
	_RegFile_reg_11__10__m2s, _RegFile_reg_11__11__m2s, _RegFile_reg_11__12__m2s,
	_RegFile_reg_11__13__m2s, _RegFile_reg_11__14__m2s, _RegFile_reg_11__15__m2s,
	_RegFile_reg_11__16__m2s, _RegFile_reg_11__17__m2s, _RegFile_reg_11__18__m2s,
	_RegFile_reg_11__19__m2s, _RegFile_reg_11__1__m2s, _RegFile_reg_11__20__m2s,
	_RegFile_reg_11__21__m2s, _RegFile_reg_11__22__m2s, _RegFile_reg_11__23__m2s,
	_RegFile_reg_11__24__m2s, _RegFile_reg_11__25__m2s, _RegFile_reg_11__26__m2s,
	_RegFile_reg_11__27__m2s, _RegFile_reg_11__28__m2s, _RegFile_reg_11__29__m2s,
	_RegFile_reg_11__2__m2s, _RegFile_reg_11__30__m2s, _RegFile_reg_11__31__m2s,
	_RegFile_reg_11__3__m2s, _RegFile_reg_11__4__m2s, _RegFile_reg_11__5__m2s,
	_RegFile_reg_11__6__m2s, _RegFile_reg_11__7__m2s, _RegFile_reg_11__8__m2s,
	_RegFile_reg_11__9__m2s, _RegFile_reg_12__0__m2s, _RegFile_reg_12__10__m2s,
	_RegFile_reg_12__11__m2s, _RegFile_reg_12__12__m2s, _RegFile_reg_12__13__m2s,
	_RegFile_reg_12__14__m2s, _RegFile_reg_12__15__m2s, _RegFile_reg_12__16__m2s,
	_RegFile_reg_12__17__m2s, _RegFile_reg_12__18__m2s, _RegFile_reg_12__19__m2s,
	_RegFile_reg_12__1__m2s, _RegFile_reg_12__20__m2s, _RegFile_reg_12__21__m2s,
	_RegFile_reg_12__22__m2s, _RegFile_reg_12__23__m2s, _RegFile_reg_12__24__m2s,
	_RegFile_reg_12__25__m2s, _RegFile_reg_12__26__m2s, _RegFile_reg_12__27__m2s,
	_RegFile_reg_12__28__m2s, _RegFile_reg_12__29__m2s, _RegFile_reg_12__2__m2s,
	_RegFile_reg_12__30__m2s, _RegFile_reg_12__31__m2s, _RegFile_reg_12__3__m2s,
	_RegFile_reg_12__4__m2s, _RegFile_reg_12__5__m2s, _RegFile_reg_12__6__m2s,
	_RegFile_reg_12__7__m2s, _RegFile_reg_12__8__m2s, _RegFile_reg_12__9__m2s,
	_RegFile_reg_13__0__m2s, _RegFile_reg_13__10__m2s, _RegFile_reg_13__11__m2s,
	_RegFile_reg_13__12__m2s, _RegFile_reg_13__13__m2s, _RegFile_reg_13__14__m2s,
	_RegFile_reg_13__15__m2s, _RegFile_reg_13__16__m2s, _RegFile_reg_13__17__m2s,
	_RegFile_reg_13__18__m2s, _RegFile_reg_13__19__m2s, _RegFile_reg_13__1__m2s,
	_RegFile_reg_13__20__m2s, _RegFile_reg_13__21__m2s, _RegFile_reg_13__22__m2s,
	_RegFile_reg_13__23__m2s, _RegFile_reg_13__24__m2s, _RegFile_reg_13__25__m2s,
	_RegFile_reg_13__26__m2s, _RegFile_reg_13__27__m2s, _RegFile_reg_13__28__m2s,
	_RegFile_reg_13__29__m2s, _RegFile_reg_13__2__m2s, _RegFile_reg_13__30__m2s,
	_RegFile_reg_13__31__m2s, _RegFile_reg_13__3__m2s, _RegFile_reg_13__4__m2s,
	_RegFile_reg_13__5__m2s, _RegFile_reg_13__6__m2s, _RegFile_reg_13__7__m2s,
	_RegFile_reg_13__8__m2s, _RegFile_reg_13__9__m2s, _RegFile_reg_14__0__m2s,
	_RegFile_reg_14__10__m2s, _RegFile_reg_14__11__m2s, _RegFile_reg_14__12__m2s,
	_RegFile_reg_14__13__m2s, _RegFile_reg_14__14__m2s, _RegFile_reg_14__15__m2s,
	_RegFile_reg_14__16__m2s, _RegFile_reg_14__17__m2s, _RegFile_reg_14__18__m2s,
	_RegFile_reg_14__19__m2s, _RegFile_reg_14__1__m2s, _RegFile_reg_14__20__m2s,
	_RegFile_reg_14__21__m2s, _RegFile_reg_14__22__m2s, _RegFile_reg_14__23__m2s,
	_RegFile_reg_14__24__m2s, _RegFile_reg_14__25__m2s, _RegFile_reg_14__26__m2s,
	_RegFile_reg_14__27__m2s, _RegFile_reg_14__28__m2s, _RegFile_reg_14__29__m2s,
	_RegFile_reg_14__2__m2s, _RegFile_reg_14__30__m2s, _RegFile_reg_14__31__m2s,
	_RegFile_reg_14__3__m2s, _RegFile_reg_14__4__m2s, _RegFile_reg_14__5__m2s,
	_RegFile_reg_14__6__m2s, _RegFile_reg_14__7__m2s, _RegFile_reg_14__8__m2s,
	_RegFile_reg_14__9__m2s, _RegFile_reg_15__0__m2s, _RegFile_reg_15__10__m2s,
	_RegFile_reg_15__11__m2s, _RegFile_reg_15__12__m2s, _RegFile_reg_15__13__m2s,
	_RegFile_reg_15__14__m2s, _RegFile_reg_15__15__m2s, _RegFile_reg_15__16__m2s,
	_RegFile_reg_15__17__m2s, _RegFile_reg_15__18__m2s, _RegFile_reg_15__19__m2s,
	_RegFile_reg_15__1__m2s, _RegFile_reg_15__20__m2s, _RegFile_reg_15__21__m2s,
	_RegFile_reg_15__22__m2s, _RegFile_reg_15__23__m2s, _RegFile_reg_15__24__m2s,
	_RegFile_reg_15__25__m2s, _RegFile_reg_15__26__m2s, _RegFile_reg_15__27__m2s,
	_RegFile_reg_15__28__m2s, _RegFile_reg_15__29__m2s, _RegFile_reg_15__2__m2s,
	_RegFile_reg_15__30__m2s, _RegFile_reg_15__31__m2s, _RegFile_reg_15__3__m2s,
	_RegFile_reg_15__4__m2s, _RegFile_reg_15__5__m2s, _RegFile_reg_15__6__m2s,
	_RegFile_reg_15__7__m2s, _RegFile_reg_15__8__m2s, _RegFile_reg_15__9__m2s,
	_RegFile_reg_16__0__m2s, _RegFile_reg_16__10__m2s, _RegFile_reg_16__11__m2s,
	_RegFile_reg_16__12__m2s, _RegFile_reg_16__13__m2s, _RegFile_reg_16__14__m2s,
	_RegFile_reg_16__15__m2s, _RegFile_reg_16__16__m2s, _RegFile_reg_16__17__m2s,
	_RegFile_reg_16__18__m2s, _RegFile_reg_16__19__m2s, _RegFile_reg_16__1__m2s,
	_RegFile_reg_16__20__m2s, _RegFile_reg_16__21__m2s, _RegFile_reg_16__22__m2s,
	_RegFile_reg_16__23__m2s, _RegFile_reg_16__24__m2s, _RegFile_reg_16__25__m2s,
	_RegFile_reg_16__26__m2s, _RegFile_reg_16__27__m2s, _RegFile_reg_16__28__m2s,
	_RegFile_reg_16__29__m2s, _RegFile_reg_16__2__m2s, _RegFile_reg_16__30__m2s,
	_RegFile_reg_16__31__m2s, _RegFile_reg_16__3__m2s, _RegFile_reg_16__4__m2s,
	_RegFile_reg_16__5__m2s, _RegFile_reg_16__6__m2s, _RegFile_reg_16__7__m2s,
	_RegFile_reg_16__8__m2s, _RegFile_reg_16__9__m2s, _RegFile_reg_17__0__m2s,
	_RegFile_reg_17__10__m2s, _RegFile_reg_17__11__m2s, _RegFile_reg_17__12__m2s,
	_RegFile_reg_17__13__m2s, _RegFile_reg_17__14__m2s, _RegFile_reg_17__15__m2s,
	_RegFile_reg_17__16__m2s, _RegFile_reg_17__17__m2s, _RegFile_reg_17__18__m2s,
	_RegFile_reg_17__19__m2s, _RegFile_reg_17__1__m2s, _RegFile_reg_17__20__m2s,
	_RegFile_reg_17__21__m2s, _RegFile_reg_17__22__m2s, _RegFile_reg_17__23__m2s,
	_RegFile_reg_17__24__m2s, _RegFile_reg_17__25__m2s, _RegFile_reg_17__26__m2s,
	_RegFile_reg_17__27__m2s, _RegFile_reg_17__28__m2s, _RegFile_reg_17__29__m2s,
	_RegFile_reg_17__2__m2s, _RegFile_reg_17__30__m2s, _RegFile_reg_17__31__m2s,
	_RegFile_reg_17__3__m2s, _RegFile_reg_17__4__m2s, _RegFile_reg_17__5__m2s,
	_RegFile_reg_17__6__m2s, _RegFile_reg_17__7__m2s, _RegFile_reg_17__8__m2s,
	_RegFile_reg_17__9__m2s, _RegFile_reg_18__0__m2s, _RegFile_reg_18__10__m2s,
	_RegFile_reg_18__11__m2s, _RegFile_reg_18__12__m2s, _RegFile_reg_18__13__m2s,
	_RegFile_reg_18__14__m2s, _RegFile_reg_18__15__m2s, _RegFile_reg_18__16__m2s,
	_RegFile_reg_18__17__m2s, _RegFile_reg_18__18__m2s, _RegFile_reg_18__19__m2s,
	_RegFile_reg_18__1__m2s, _RegFile_reg_18__20__m2s, _RegFile_reg_18__21__m2s,
	_RegFile_reg_18__22__m2s, _RegFile_reg_18__23__m2s, _RegFile_reg_18__24__m2s,
	_RegFile_reg_18__25__m2s, _RegFile_reg_18__26__m2s, _RegFile_reg_18__27__m2s,
	_RegFile_reg_18__28__m2s, _RegFile_reg_18__29__m2s, _RegFile_reg_18__2__m2s,
	_RegFile_reg_18__30__m2s, _RegFile_reg_18__31__m2s, _RegFile_reg_18__3__m2s,
	_RegFile_reg_18__4__m2s, _RegFile_reg_18__5__m2s, _RegFile_reg_18__6__m2s,
	_RegFile_reg_18__7__m2s, _RegFile_reg_18__8__m2s, _RegFile_reg_18__9__m2s,
	_RegFile_reg_19__0__m2s, _RegFile_reg_19__10__m2s, _RegFile_reg_19__11__m2s,
	_RegFile_reg_19__12__m2s, _RegFile_reg_19__13__m2s, _RegFile_reg_19__14__m2s,
	_RegFile_reg_19__15__m2s, _RegFile_reg_19__16__m2s, _RegFile_reg_19__17__m2s,
	_RegFile_reg_19__18__m2s, _RegFile_reg_19__19__m2s, _RegFile_reg_19__1__m2s,
	_RegFile_reg_19__20__m2s, _RegFile_reg_19__21__m2s, _RegFile_reg_19__22__m2s,
	_RegFile_reg_19__23__m2s, _RegFile_reg_19__24__m2s, _RegFile_reg_19__25__m2s,
	_RegFile_reg_19__26__m2s, _RegFile_reg_19__27__m2s, _RegFile_reg_19__28__m2s,
	_RegFile_reg_19__29__m2s, _RegFile_reg_19__2__m2s, _RegFile_reg_19__30__m2s,
	_RegFile_reg_19__31__m2s, _RegFile_reg_19__3__m2s, _RegFile_reg_19__4__m2s,
	_RegFile_reg_19__5__m2s, _RegFile_reg_19__6__m2s, _RegFile_reg_19__7__m2s,
	_RegFile_reg_19__8__m2s, _RegFile_reg_19__9__m2s, _RegFile_reg_1__0__m2s,
	_RegFile_reg_1__10__m2s, _RegFile_reg_1__11__m2s, _RegFile_reg_1__12__m2s,
	_RegFile_reg_1__13__m2s, _RegFile_reg_1__14__m2s, _RegFile_reg_1__15__m2s,
	_RegFile_reg_1__16__m2s, _RegFile_reg_1__17__m2s, _RegFile_reg_1__18__m2s,
	_RegFile_reg_1__19__m2s, _RegFile_reg_1__1__m2s, _RegFile_reg_1__20__m2s,
	_RegFile_reg_1__21__m2s, _RegFile_reg_1__22__m2s, _RegFile_reg_1__23__m2s,
	_RegFile_reg_1__24__m2s, _RegFile_reg_1__25__m2s, _RegFile_reg_1__26__m2s,
	_RegFile_reg_1__27__m2s, _RegFile_reg_1__28__m2s, _RegFile_reg_1__29__m2s,
	_RegFile_reg_1__2__m2s, _RegFile_reg_1__30__m2s, _RegFile_reg_1__31__m2s,
	_RegFile_reg_1__3__m2s, _RegFile_reg_1__4__m2s, _RegFile_reg_1__5__m2s,
	_RegFile_reg_1__6__m2s, _RegFile_reg_1__7__m2s, _RegFile_reg_1__8__m2s,
	_RegFile_reg_1__9__m2s, _RegFile_reg_20__0__m2s, _RegFile_reg_20__10__m2s,
	_RegFile_reg_20__11__m2s, _RegFile_reg_20__12__m2s, _RegFile_reg_20__13__m2s,
	_RegFile_reg_20__14__m2s, _RegFile_reg_20__15__m2s, _RegFile_reg_20__16__m2s,
	_RegFile_reg_20__17__m2s, _RegFile_reg_20__18__m2s, _RegFile_reg_20__19__m2s,
	_RegFile_reg_20__1__m2s, _RegFile_reg_20__20__m2s, _RegFile_reg_20__21__m2s,
	_RegFile_reg_20__22__m2s, _RegFile_reg_20__23__m2s, _RegFile_reg_20__24__m2s,
	_RegFile_reg_20__25__m2s, _RegFile_reg_20__26__m2s, _RegFile_reg_20__27__m2s,
	_RegFile_reg_20__28__m2s, _RegFile_reg_20__29__m2s, _RegFile_reg_20__2__m2s,
	_RegFile_reg_20__30__m2s, _RegFile_reg_20__31__m2s, _RegFile_reg_20__3__m2s,
	_RegFile_reg_20__4__m2s, _RegFile_reg_20__5__m2s, _RegFile_reg_20__6__m2s,
	_RegFile_reg_20__7__m2s, _RegFile_reg_20__8__m2s, _RegFile_reg_20__9__m2s,
	_RegFile_reg_21__0__m2s, _RegFile_reg_21__10__m2s, _RegFile_reg_21__11__m2s,
	_RegFile_reg_21__12__m2s, _RegFile_reg_21__13__m2s, _RegFile_reg_21__14__m2s,
	_RegFile_reg_21__15__m2s, _RegFile_reg_21__16__m2s, _RegFile_reg_21__17__m2s,
	_RegFile_reg_21__18__m2s, _RegFile_reg_21__19__m2s, _RegFile_reg_21__1__m2s,
	_RegFile_reg_21__20__m2s, _RegFile_reg_21__21__m2s, _RegFile_reg_21__22__m2s,
	_RegFile_reg_21__23__m2s, _RegFile_reg_21__24__m2s, _RegFile_reg_21__25__m2s,
	_RegFile_reg_21__26__m2s, _RegFile_reg_21__27__m2s, _RegFile_reg_21__28__m2s,
	_RegFile_reg_21__29__m2s, _RegFile_reg_21__2__m2s, _RegFile_reg_21__30__m2s,
	_RegFile_reg_21__31__m2s, _RegFile_reg_21__3__m2s, _RegFile_reg_21__4__m2s,
	_RegFile_reg_21__5__m2s, _RegFile_reg_21__6__m2s, _RegFile_reg_21__7__m2s,
	_RegFile_reg_21__8__m2s, _RegFile_reg_21__9__m2s, _RegFile_reg_22__0__m2s,
	_RegFile_reg_22__10__m2s, _RegFile_reg_22__11__m2s, _RegFile_reg_22__12__m2s,
	_RegFile_reg_22__13__m2s, _RegFile_reg_22__14__m2s, _RegFile_reg_22__15__m2s,
	_RegFile_reg_22__16__m2s, _RegFile_reg_22__17__m2s, _RegFile_reg_22__18__m2s,
	_RegFile_reg_22__19__m2s, _RegFile_reg_22__1__m2s, _RegFile_reg_22__20__m2s,
	_RegFile_reg_22__21__m2s, _RegFile_reg_22__22__m2s, _RegFile_reg_22__23__m2s,
	_RegFile_reg_22__24__m2s, _RegFile_reg_22__25__m2s, _RegFile_reg_22__26__m2s,
	_RegFile_reg_22__27__m2s, _RegFile_reg_22__28__m2s, _RegFile_reg_22__29__m2s,
	_RegFile_reg_22__2__m2s, _RegFile_reg_22__30__m2s, _RegFile_reg_22__31__m2s,
	_RegFile_reg_22__3__m2s, _RegFile_reg_22__4__m2s, _RegFile_reg_22__5__m2s,
	_RegFile_reg_22__6__m2s, _RegFile_reg_22__7__m2s, _RegFile_reg_22__8__m2s,
	_RegFile_reg_22__9__m2s, _RegFile_reg_23__0__m2s, _RegFile_reg_23__10__m2s,
	_RegFile_reg_23__11__m2s, _RegFile_reg_23__12__m2s, _RegFile_reg_23__13__m2s,
	_RegFile_reg_23__14__m2s, _RegFile_reg_23__15__m2s, _RegFile_reg_23__16__m2s,
	_RegFile_reg_23__17__m2s, _RegFile_reg_23__18__m2s, _RegFile_reg_23__19__m2s,
	_RegFile_reg_23__1__m2s, _RegFile_reg_23__20__m2s, _RegFile_reg_23__21__m2s,
	_RegFile_reg_23__22__m2s, _RegFile_reg_23__23__m2s, _RegFile_reg_23__24__m2s,
	_RegFile_reg_23__25__m2s, _RegFile_reg_23__26__m2s, _RegFile_reg_23__27__m2s,
	_RegFile_reg_23__28__m2s, _RegFile_reg_23__29__m2s, _RegFile_reg_23__2__m2s,
	_RegFile_reg_23__30__m2s, _RegFile_reg_23__31__m2s, _RegFile_reg_23__3__m2s,
	_RegFile_reg_23__4__m2s, _RegFile_reg_23__5__m2s, _RegFile_reg_23__6__m2s,
	_RegFile_reg_23__7__m2s, _RegFile_reg_23__8__m2s, _RegFile_reg_23__9__m2s,
	_RegFile_reg_24__0__m2s, _RegFile_reg_24__10__m2s, _RegFile_reg_24__11__m2s,
	_RegFile_reg_24__12__m2s, _RegFile_reg_24__13__m2s, _RegFile_reg_24__14__m2s,
	_RegFile_reg_24__15__m2s, _RegFile_reg_24__16__m2s, _RegFile_reg_24__17__m2s,
	_RegFile_reg_24__18__m2s, _RegFile_reg_24__19__m2s, _RegFile_reg_24__1__m2s,
	_RegFile_reg_24__20__m2s, _RegFile_reg_24__21__m2s, _RegFile_reg_24__22__m2s,
	_RegFile_reg_24__23__m2s, _RegFile_reg_24__24__m2s, _RegFile_reg_24__25__m2s,
	_RegFile_reg_24__26__m2s, _RegFile_reg_24__27__m2s, _RegFile_reg_24__28__m2s,
	_RegFile_reg_24__29__m2s, _RegFile_reg_24__2__m2s, _RegFile_reg_24__30__m2s,
	_RegFile_reg_24__31__m2s, _RegFile_reg_24__3__m2s, _RegFile_reg_24__4__m2s,
	_RegFile_reg_24__5__m2s, _RegFile_reg_24__6__m2s, _RegFile_reg_24__7__m2s,
	_RegFile_reg_24__8__m2s, _RegFile_reg_24__9__m2s, _RegFile_reg_25__0__m2s,
	_RegFile_reg_25__10__m2s, _RegFile_reg_25__11__m2s, _RegFile_reg_25__12__m2s,
	_RegFile_reg_25__13__m2s, _RegFile_reg_25__14__m2s, _RegFile_reg_25__15__m2s,
	_RegFile_reg_25__16__m2s, _RegFile_reg_25__17__m2s, _RegFile_reg_25__18__m2s,
	_RegFile_reg_25__19__m2s, _RegFile_reg_25__1__m2s, _RegFile_reg_25__20__m2s,
	_RegFile_reg_25__21__m2s, _RegFile_reg_25__22__m2s, _RegFile_reg_25__23__m2s,
	_RegFile_reg_25__24__m2s, _RegFile_reg_25__25__m2s, _RegFile_reg_25__26__m2s,
	_RegFile_reg_25__27__m2s, _RegFile_reg_25__28__m2s, _RegFile_reg_25__29__m2s,
	_RegFile_reg_25__2__m2s, _RegFile_reg_25__30__m2s, _RegFile_reg_25__31__m2s,
	_RegFile_reg_25__3__m2s, _RegFile_reg_25__4__m2s, _RegFile_reg_25__5__m2s,
	_RegFile_reg_25__6__m2s, _RegFile_reg_25__7__m2s, _RegFile_reg_25__8__m2s,
	_RegFile_reg_25__9__m2s, _RegFile_reg_26__0__m2s, _RegFile_reg_26__10__m2s,
	_RegFile_reg_26__11__m2s, _RegFile_reg_26__12__m2s, _RegFile_reg_26__13__m2s,
	_RegFile_reg_26__14__m2s, _RegFile_reg_26__15__m2s, _RegFile_reg_26__16__m2s,
	_RegFile_reg_26__17__m2s, _RegFile_reg_26__18__m2s, _RegFile_reg_26__19__m2s,
	_RegFile_reg_26__1__m2s, _RegFile_reg_26__20__m2s, _RegFile_reg_26__21__m2s,
	_RegFile_reg_26__22__m2s, _RegFile_reg_26__23__m2s, _RegFile_reg_26__24__m2s,
	_RegFile_reg_26__25__m2s, _RegFile_reg_26__26__m2s, _RegFile_reg_26__27__m2s,
	_RegFile_reg_26__28__m2s, _RegFile_reg_26__29__m2s, _RegFile_reg_26__2__m2s,
	_RegFile_reg_26__30__m2s, _RegFile_reg_26__31__m2s, _RegFile_reg_26__3__m2s,
	_RegFile_reg_26__4__m2s, _RegFile_reg_26__5__m2s, _RegFile_reg_26__6__m2s,
	_RegFile_reg_26__7__m2s, _RegFile_reg_26__8__m2s, _RegFile_reg_26__9__m2s,
	_RegFile_reg_27__0__m2s, _RegFile_reg_27__10__m2s, _RegFile_reg_27__11__m2s,
	_RegFile_reg_27__12__m2s, _RegFile_reg_27__13__m2s, _RegFile_reg_27__14__m2s,
	_RegFile_reg_27__15__m2s, _RegFile_reg_27__16__m2s, _RegFile_reg_27__17__m2s,
	_RegFile_reg_27__18__m2s, _RegFile_reg_27__19__m2s, _RegFile_reg_27__1__m2s,
	_RegFile_reg_27__20__m2s, _RegFile_reg_27__21__m2s, _RegFile_reg_27__22__m2s,
	_RegFile_reg_27__23__m2s, _RegFile_reg_27__24__m2s, _RegFile_reg_27__25__m2s,
	_RegFile_reg_27__26__m2s, _RegFile_reg_27__27__m2s, _RegFile_reg_27__28__m2s,
	_RegFile_reg_27__29__m2s, _RegFile_reg_27__2__m2s, _RegFile_reg_27__30__m2s,
	_RegFile_reg_27__31__m2s, _RegFile_reg_27__3__m2s, _RegFile_reg_27__4__m2s,
	_RegFile_reg_27__5__m2s, _RegFile_reg_27__6__m2s, _RegFile_reg_27__7__m2s,
	_RegFile_reg_27__8__m2s, _RegFile_reg_27__9__m2s, _RegFile_reg_28__0__m2s,
	_RegFile_reg_28__10__m2s, _RegFile_reg_28__11__m2s, _RegFile_reg_28__12__m2s,
	_RegFile_reg_28__13__m2s, _RegFile_reg_28__14__m2s, _RegFile_reg_28__15__m2s,
	_RegFile_reg_28__16__m2s, _RegFile_reg_28__17__m2s, _RegFile_reg_28__18__m2s,
	_RegFile_reg_28__19__m2s, _RegFile_reg_28__1__m2s, _RegFile_reg_28__20__m2s,
	_RegFile_reg_28__21__m2s, _RegFile_reg_28__22__m2s, _RegFile_reg_28__23__m2s,
	_RegFile_reg_28__24__m2s, _RegFile_reg_28__25__m2s, _RegFile_reg_28__26__m2s,
	_RegFile_reg_28__27__m2s, _RegFile_reg_28__28__m2s, _RegFile_reg_28__29__m2s,
	_RegFile_reg_28__2__m2s, _RegFile_reg_28__30__m2s, _RegFile_reg_28__31__m2s,
	_RegFile_reg_28__3__m2s, _RegFile_reg_28__4__m2s, _RegFile_reg_28__5__m2s,
	_RegFile_reg_28__6__m2s, _RegFile_reg_28__7__m2s, _RegFile_reg_28__8__m2s,
	_RegFile_reg_28__9__m2s, _RegFile_reg_29__0__m2s, _RegFile_reg_29__10__m2s,
	_RegFile_reg_29__11__m2s, _RegFile_reg_29__12__m2s, _RegFile_reg_29__13__m2s,
	_RegFile_reg_29__14__m2s, _RegFile_reg_29__15__m2s, _RegFile_reg_29__16__m2s,
	_RegFile_reg_29__17__m2s, _RegFile_reg_29__18__m2s, _RegFile_reg_29__19__m2s,
	_RegFile_reg_29__1__m2s, _RegFile_reg_29__20__m2s, _RegFile_reg_29__21__m2s,
	_RegFile_reg_29__22__m2s, _RegFile_reg_29__23__m2s, _RegFile_reg_29__24__m2s,
	_RegFile_reg_29__25__m2s, _RegFile_reg_29__26__m2s, _RegFile_reg_29__27__m2s,
	_RegFile_reg_29__28__m2s, _RegFile_reg_29__29__m2s, _RegFile_reg_29__2__m2s,
	_RegFile_reg_29__30__m2s, _RegFile_reg_29__31__m2s, _RegFile_reg_29__3__m2s,
	_RegFile_reg_29__4__m2s, _RegFile_reg_29__5__m2s, _RegFile_reg_29__6__m2s,
	_RegFile_reg_29__7__m2s, _RegFile_reg_29__8__m2s, _RegFile_reg_29__9__m2s,
	_RegFile_reg_2__0__m2s, _RegFile_reg_2__10__m2s, _RegFile_reg_2__11__m2s,
	_RegFile_reg_2__12__m2s, _RegFile_reg_2__13__m2s, _RegFile_reg_2__14__m2s,
	_RegFile_reg_2__15__m2s, _RegFile_reg_2__16__m2s, _RegFile_reg_2__17__m2s,
	_RegFile_reg_2__18__m2s, _RegFile_reg_2__19__m2s, _RegFile_reg_2__1__m2s,
	_RegFile_reg_2__20__m2s, _RegFile_reg_2__21__m2s, _RegFile_reg_2__22__m2s,
	_RegFile_reg_2__23__m2s, _RegFile_reg_2__24__m2s, _RegFile_reg_2__25__m2s,
	_RegFile_reg_2__26__m2s, _RegFile_reg_2__27__m2s, _RegFile_reg_2__28__m2s,
	_RegFile_reg_2__29__m2s, _RegFile_reg_2__2__m2s, _RegFile_reg_2__30__m2s,
	_RegFile_reg_2__31__m2s, _RegFile_reg_2__3__m2s, _RegFile_reg_2__4__m2s,
	_RegFile_reg_2__5__m2s, _RegFile_reg_2__6__m2s, _RegFile_reg_2__7__m2s,
	_RegFile_reg_2__8__m2s, _RegFile_reg_2__9__m2s, _RegFile_reg_30__0__m2s,
	_RegFile_reg_30__10__m2s, _RegFile_reg_30__11__m2s, _RegFile_reg_30__12__m2s,
	_RegFile_reg_30__13__m2s, _RegFile_reg_30__14__m2s, _RegFile_reg_30__15__m2s,
	_RegFile_reg_30__16__m2s, _RegFile_reg_30__17__m2s, _RegFile_reg_30__18__m2s,
	_RegFile_reg_30__19__m2s, _RegFile_reg_30__1__m2s, _RegFile_reg_30__20__m2s,
	_RegFile_reg_30__21__m2s, _RegFile_reg_30__22__m2s, _RegFile_reg_30__23__m2s,
	_RegFile_reg_30__24__m2s, _RegFile_reg_30__25__m2s, _RegFile_reg_30__26__m2s,
	_RegFile_reg_30__27__m2s, _RegFile_reg_30__28__m2s, _RegFile_reg_30__29__m2s,
	_RegFile_reg_30__2__m2s, _RegFile_reg_30__30__m2s, _RegFile_reg_30__31__m2s,
	_RegFile_reg_30__3__m2s, _RegFile_reg_30__4__m2s, _RegFile_reg_30__5__m2s,
	_RegFile_reg_30__6__m2s, _RegFile_reg_30__7__m2s, _RegFile_reg_30__8__m2s,
	_RegFile_reg_30__9__m2s, _RegFile_reg_31__0__m2s, _RegFile_reg_31__10__m2s,
	_RegFile_reg_31__11__m2s, _RegFile_reg_31__12__m2s, _RegFile_reg_31__13__m2s,
	_RegFile_reg_31__14__m2s, _RegFile_reg_31__15__m2s, _RegFile_reg_31__16__m2s,
	_RegFile_reg_31__17__m2s, _RegFile_reg_31__18__m2s, _RegFile_reg_31__19__m2s,
	_RegFile_reg_31__1__m2s, _RegFile_reg_31__20__m2s, _RegFile_reg_31__21__m2s,
	_RegFile_reg_31__22__m2s, _RegFile_reg_31__23__m2s, _RegFile_reg_31__24__m2s,
	_RegFile_reg_31__25__m2s, _RegFile_reg_31__26__m2s, _RegFile_reg_31__27__m2s,
	_RegFile_reg_31__28__m2s, _RegFile_reg_31__29__m2s, _RegFile_reg_31__2__m2s,
	_RegFile_reg_31__30__m2s, _RegFile_reg_31__31__m2s, _RegFile_reg_31__3__m2s,
	_RegFile_reg_31__4__m2s, _RegFile_reg_31__5__m2s, _RegFile_reg_31__6__m2s,
	_RegFile_reg_31__7__m2s, _RegFile_reg_31__8__m2s, _RegFile_reg_31__9__m2s,
	_RegFile_reg_3__0__m2s, _RegFile_reg_3__10__m2s, _RegFile_reg_3__11__m2s,
	_RegFile_reg_3__12__m2s, _RegFile_reg_3__13__m2s, _RegFile_reg_3__14__m2s,
	_RegFile_reg_3__15__m2s, _RegFile_reg_3__16__m2s, _RegFile_reg_3__17__m2s,
	_RegFile_reg_3__18__m2s, _RegFile_reg_3__19__m2s, _RegFile_reg_3__1__m2s,
	_RegFile_reg_3__20__m2s, _RegFile_reg_3__21__m2s, _RegFile_reg_3__22__m2s,
	_RegFile_reg_3__23__m2s, _RegFile_reg_3__24__m2s, _RegFile_reg_3__25__m2s,
	_RegFile_reg_3__26__m2s, _RegFile_reg_3__27__m2s, _RegFile_reg_3__28__m2s,
	_RegFile_reg_3__29__m2s, _RegFile_reg_3__2__m2s, _RegFile_reg_3__30__m2s,
	_RegFile_reg_3__31__m2s, _RegFile_reg_3__3__m2s, _RegFile_reg_3__4__m2s,
	_RegFile_reg_3__5__m2s, _RegFile_reg_3__6__m2s, _RegFile_reg_3__7__m2s,
	_RegFile_reg_3__8__m2s, _RegFile_reg_3__9__m2s, _RegFile_reg_4__0__m2s,
	_RegFile_reg_4__10__m2s, _RegFile_reg_4__11__m2s, _RegFile_reg_4__12__m2s,
	_RegFile_reg_4__13__m2s, _RegFile_reg_4__14__m2s, _RegFile_reg_4__15__m2s,
	_RegFile_reg_4__16__m2s, _RegFile_reg_4__17__m2s, _RegFile_reg_4__18__m2s,
	_RegFile_reg_4__19__m2s, _RegFile_reg_4__1__m2s, _RegFile_reg_4__20__m2s,
	_RegFile_reg_4__21__m2s, _RegFile_reg_4__22__m2s, _RegFile_reg_4__23__m2s,
	_RegFile_reg_4__24__m2s, _RegFile_reg_4__25__m2s, _RegFile_reg_4__26__m2s,
	_RegFile_reg_4__27__m2s, _RegFile_reg_4__28__m2s, _RegFile_reg_4__29__m2s,
	_RegFile_reg_4__2__m2s, _RegFile_reg_4__30__m2s, _RegFile_reg_4__31__m2s,
	_RegFile_reg_4__3__m2s, _RegFile_reg_4__4__m2s, _RegFile_reg_4__5__m2s,
	_RegFile_reg_4__6__m2s, _RegFile_reg_4__7__m2s, _RegFile_reg_4__8__m2s,
	_RegFile_reg_4__9__m2s, _RegFile_reg_5__0__m2s, _RegFile_reg_5__10__m2s,
	_RegFile_reg_5__11__m2s, _RegFile_reg_5__12__m2s, _RegFile_reg_5__13__m2s,
	_RegFile_reg_5__14__m2s, _RegFile_reg_5__15__m2s, _RegFile_reg_5__16__m2s,
	_RegFile_reg_5__17__m2s, _RegFile_reg_5__18__m2s, _RegFile_reg_5__19__m2s,
	_RegFile_reg_5__1__m2s, _RegFile_reg_5__20__m2s, _RegFile_reg_5__21__m2s,
	_RegFile_reg_5__22__m2s, _RegFile_reg_5__23__m2s, _RegFile_reg_5__24__m2s,
	_RegFile_reg_5__25__m2s, _RegFile_reg_5__26__m2s, _RegFile_reg_5__27__m2s,
	_RegFile_reg_5__28__m2s, _RegFile_reg_5__29__m2s, _RegFile_reg_5__2__m2s,
	_RegFile_reg_5__30__m2s, _RegFile_reg_5__31__m2s, _RegFile_reg_5__3__m2s,
	_RegFile_reg_5__4__m2s, _RegFile_reg_5__5__m2s, _RegFile_reg_5__6__m2s,
	_RegFile_reg_5__7__m2s, _RegFile_reg_5__8__m2s, _RegFile_reg_5__9__m2s,
	_RegFile_reg_6__0__m2s, _RegFile_reg_6__10__m2s, _RegFile_reg_6__11__m2s,
	_RegFile_reg_6__12__m2s, _RegFile_reg_6__13__m2s, _RegFile_reg_6__14__m2s,
	_RegFile_reg_6__15__m2s, _RegFile_reg_6__16__m2s, _RegFile_reg_6__17__m2s,
	_RegFile_reg_6__18__m2s, _RegFile_reg_6__19__m2s, _RegFile_reg_6__1__m2s,
	_RegFile_reg_6__20__m2s, _RegFile_reg_6__21__m2s, _RegFile_reg_6__22__m2s,
	_RegFile_reg_6__23__m2s, _RegFile_reg_6__24__m2s, _RegFile_reg_6__25__m2s,
	_RegFile_reg_6__26__m2s, _RegFile_reg_6__27__m2s, _RegFile_reg_6__28__m2s,
	_RegFile_reg_6__29__m2s, _RegFile_reg_6__2__m2s, _RegFile_reg_6__30__m2s,
	_RegFile_reg_6__31__m2s, _RegFile_reg_6__3__m2s, _RegFile_reg_6__4__m2s,
	_RegFile_reg_6__5__m2s, _RegFile_reg_6__6__m2s, _RegFile_reg_6__7__m2s,
	_RegFile_reg_6__8__m2s, _RegFile_reg_6__9__m2s, _RegFile_reg_7__0__m2s,
	_RegFile_reg_7__10__m2s, _RegFile_reg_7__11__m2s, _RegFile_reg_7__12__m2s,
	_RegFile_reg_7__13__m2s, _RegFile_reg_7__14__m2s, _RegFile_reg_7__15__m2s,
	_RegFile_reg_7__16__m2s, _RegFile_reg_7__17__m2s, _RegFile_reg_7__18__m2s,
	_RegFile_reg_7__19__m2s, _RegFile_reg_7__1__m2s, _RegFile_reg_7__20__m2s,
	_RegFile_reg_7__21__m2s, _RegFile_reg_7__22__m2s, _RegFile_reg_7__23__m2s,
	_RegFile_reg_7__24__m2s, _RegFile_reg_7__25__m2s, _RegFile_reg_7__26__m2s,
	_RegFile_reg_7__27__m2s, _RegFile_reg_7__28__m2s, _RegFile_reg_7__29__m2s,
	_RegFile_reg_7__2__m2s, _RegFile_reg_7__30__m2s, _RegFile_reg_7__31__m2s,
	_RegFile_reg_7__3__m2s, _RegFile_reg_7__4__m2s, _RegFile_reg_7__5__m2s,
	_RegFile_reg_7__6__m2s, _RegFile_reg_7__7__m2s, _RegFile_reg_7__8__m2s,
	_RegFile_reg_7__9__m2s, _RegFile_reg_8__0__m2s, _RegFile_reg_8__10__m2s,
	_RegFile_reg_8__11__m2s, _RegFile_reg_8__12__m2s, _RegFile_reg_8__13__m2s,
	_RegFile_reg_8__14__m2s, _RegFile_reg_8__15__m2s, _RegFile_reg_8__16__m2s,
	_RegFile_reg_8__17__m2s, _RegFile_reg_8__18__m2s, _RegFile_reg_8__19__m2s,
	_RegFile_reg_8__1__m2s, _RegFile_reg_8__20__m2s, _RegFile_reg_8__21__m2s,
	_RegFile_reg_8__22__m2s, _RegFile_reg_8__23__m2s, _RegFile_reg_8__24__m2s,
	_RegFile_reg_8__25__m2s, _RegFile_reg_8__26__m2s, _RegFile_reg_8__27__m2s,
	_RegFile_reg_8__28__m2s, _RegFile_reg_8__29__m2s, _RegFile_reg_8__2__m2s,
	_RegFile_reg_8__30__m2s, _RegFile_reg_8__31__m2s, _RegFile_reg_8__3__m2s,
	_RegFile_reg_8__4__m2s, _RegFile_reg_8__5__m2s, _RegFile_reg_8__6__m2s,
	_RegFile_reg_8__7__m2s, _RegFile_reg_8__8__m2s, _RegFile_reg_8__9__m2s,
	_RegFile_reg_9__0__m2s, _RegFile_reg_9__10__m2s, _RegFile_reg_9__11__m2s,
	_RegFile_reg_9__12__m2s, _RegFile_reg_9__13__m2s, _RegFile_reg_9__14__m2s,
	_RegFile_reg_9__15__m2s, _RegFile_reg_9__16__m2s, _RegFile_reg_9__17__m2s,
	_RegFile_reg_9__18__m2s, _RegFile_reg_9__19__m2s, _RegFile_reg_9__1__m2s,
	_RegFile_reg_9__20__m2s, _RegFile_reg_9__21__m2s, _RegFile_reg_9__22__m2s,
	_RegFile_reg_9__23__m2s, _RegFile_reg_9__24__m2s, _RegFile_reg_9__25__m2s,
	_RegFile_reg_9__26__m2s, _RegFile_reg_9__27__m2s, _RegFile_reg_9__28__m2s,
	_RegFile_reg_9__29__m2s, _RegFile_reg_9__2__m2s, _RegFile_reg_9__30__m2s,
	_RegFile_reg_9__31__m2s, _RegFile_reg_9__3__m2s, _RegFile_reg_9__4__m2s,
	_RegFile_reg_9__5__m2s, _RegFile_reg_9__6__m2s, _RegFile_reg_9__7__m2s,
	_RegFile_reg_9__8__m2s, _RegFile_reg_9__9__m2s, ___cell__36997_net125928,
	___cell__36997_net125941, ___cell__36997_net125989, ___cell__36997_net126005,
	___cell__36997_net126604, ___cell__36997_net126612, ___cell__36997_net126621,
	___cell__36997_net127155, ___cell__36997_net127189, ___cell__36997_net127190,
	___cell__36997_net127210, ___cell__36997_net129239, ___cell__36997_net129247,
	___cell__36997_net129354, ___cell__36997_net129378, ___cell__36997_net129381,
	___cell__36997_net129384, ___cell__36997_net129388, ___cell__36997_net129389,
	___cell__36997_net129477, ___cell__36997_net129524, ___cell__36997_net129624,
	___cell__36997_net129625, ___cell__36997_net129626, ___cell__36997_net129632,
	___cell__36997_net129654, ___cell__36997_net129657, ___cell__36997_net129786,
	___cell__36997_net129977, ___cell__36997_net129979, ___cell__36997_net130125,
	___cell__36997_net130187, ___cell__36997_net130191, ___cell__36997_net130212,
	___cell__36997_net130214, ___cell__36997_net130217, ___cell__36997_net130306,
	___cell__36997_net130567, ___cell__36997_net130572, ___cell__36997_net130580,
	___cell__36997_net130681, ___cell__36997_net130705, ___cell__36997_net130709,
	___cell__36997_net130713, ___cell__6171_net27367, _branch_address_reg_31_net46811,
	_counter_reg_0_net48671, _counter_reg_1_net48651, _current_IR_reg_1_net49291,
	branch_address_reg_0__m2s, branch_address_reg_10__m2s, branch_address_reg_11__m2s,
	branch_address_reg_12__m2s, branch_address_reg_13__m2s, branch_address_reg_14__m2s,
	branch_address_reg_15__m2s, branch_address_reg_16__m2s, branch_address_reg_17__m2s,
	branch_address_reg_18__m2s, branch_address_reg_19__m2s, branch_address_reg_1__m2s,
	branch_address_reg_20__m2s, branch_address_reg_21__m2s, branch_address_reg_22__m2s,
	branch_address_reg_23__m2s, branch_address_reg_24__m2s, branch_address_reg_25__m2s,
	branch_address_reg_26__m2s, branch_address_reg_27__m2s, branch_address_reg_28__m2s,
	branch_address_reg_29__m2s, branch_address_reg_2__m2s, branch_address_reg_30__m2s,
	branch_address_reg_31__m2s, branch_address_reg_3__m2s, branch_address_reg_4__m2s,
	branch_address_reg_5__m2s, branch_address_reg_6__m2s, branch_address_reg_7__m2s,
	branch_address_reg_8__m2s, branch_address_reg_9__m2s, branch_sig_reg__m2s,
	counter_reg_0__m2s, counter_reg_1__m2s, current_IR_0, current_IR_1, current_IR_10,
	current_IR_17, current_IR_18, current_IR_19, current_IR_2, current_IR_21,
	current_IR_23, current_IR_24, current_IR_27, current_IR_29, current_IR_3,
	current_IR_30, current_IR_31, current_IR_4, current_IR_6, current_IR_7,
	current_IR_8, current_IR_9, current_IR_reg_0__m2s, current_IR_reg_10__m2s,
	current_IR_reg_11__m2s, current_IR_reg_12__m2s, current_IR_reg_13__m2s,
	current_IR_reg_14__m2s, current_IR_reg_15__m2s, current_IR_reg_16__m2s,
	current_IR_reg_17__m2s, current_IR_reg_18__m2s, current_IR_reg_19__m2s,
	current_IR_reg_1__m2s, current_IR_reg_20__m2s, current_IR_reg_21__m2s,
	current_IR_reg_22__m2s, current_IR_reg_23__m2s, current_IR_reg_24__m2s,
	current_IR_reg_25__m2s, current_IR_reg_26__m2s, current_IR_reg_27__m2s,
	current_IR_reg_28__m2s, current_IR_reg_29__m2s, current_IR_reg_2__m2s,
	current_IR_reg_30__m2s, current_IR_reg_31__m2s, current_IR_reg_3__m2s,
	current_IR_reg_4__m2s, current_IR_reg_5__m2s, current_IR_reg_6__m2s, current_IR_reg_7__m2s,
	current_IR_reg_8__m2s, current_IR_reg_9__m2s, delay_slot, delay_slot_reg__m2s,
	intr_slot, intr_slot_reg__m2s, mem_read_reg__m2s, mem_to_reg_reg__m2s,
	mem_write_reg__m2s, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
	n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
	n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
	n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
	n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
	n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
	n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
	n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
	n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
	n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
	n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
	n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
	n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
	n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
	n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
	n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
	n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
	n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
	n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
	n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
	n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
	n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
	n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
	n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
	n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
	n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
	n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
	n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
	n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
	n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
	n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
	n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
	n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
	n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
	n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
	n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
	n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
	n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
	n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
	n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
	n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
	n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
	n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
	n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
	n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
	n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
	n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
	n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
	n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
	n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
	n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
	n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
	n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
	n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
	n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
	n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1557, n1558, n1559,
	n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
	n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1578, n1579, n1580,
	n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
	n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
	n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
	n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
	n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
	n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
	n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
	n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
	n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
	n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
	n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
	n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
	n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
	n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
	n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
	n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
	n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
	n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
	n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
	n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
	n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
	n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
	n1801, n1802, n1803, n1804, n1826, n1827, n1828, n1829, n1830, n1831,
	n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
	n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
	n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
	n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
	n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
	n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
	n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
	n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
	n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
	n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
	n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
	n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
	n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
	n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
	n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
	n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
	n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
	n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
	n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
	n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
	n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
	n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
	n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
	n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
	n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
	n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
	n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
	n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
	n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
	n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
	n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
	n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
	n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
	n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
	n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
	n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
	n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
	n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
	n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
	n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
	n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
	n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
	n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
	n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
	n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
	n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
	n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
	n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
	n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
	n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
	n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
	n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
	n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
	n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
	n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
	n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
	n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
	n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
	n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
	n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
	n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
	n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
	n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
	n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
	n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
	n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
	n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
	n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
	n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
	n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
	n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
	n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
	n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
	n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
	n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
	n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
	n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
	n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
	n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
	n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
	n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
	n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
	n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
	n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
	n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
	n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
	n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
	n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
	n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
	n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
	n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
	n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
	n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
	n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
	n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
	n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
	n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
	n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
	n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
	n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
	n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
	n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
	n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
	n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
	n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
	n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
	n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
	n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
	n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
	n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
	n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
	n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
	n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
	n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
	n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
	n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
	n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
	n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
	n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
	n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
	n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
	n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
	n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
	n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
	n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
	n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
	n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
	n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
	n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
	n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
	n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
	n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
	n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
	n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
	n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
	n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
	n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
	n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
	n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
	n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
	n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
	n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
	n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
	n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
	n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
	n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
	n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
	n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n331, n3310, n3311,
	n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n332, n3320, n3321,
	n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n333, n3330, n3331,
	n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n334, n3340, n3341,
	n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n335, n3350, n3351,
	n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n336, n3360, n3361,
	n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n337, n3370, n3371,
	n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n338, n3380, n3381,
	n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n339, n3390, n3391,
	n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n340, n3400, n3401,
	n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
	n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
	n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
	n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
	n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
	n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
	n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
	n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
	n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
	n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
	n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
	n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
	n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
	n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
	n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
	n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
	n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
	n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
	n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
	n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
	n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
	n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
	n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
	n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
	n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
	n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
	n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
	n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
	n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
	n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
	n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
	n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
	n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
	n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
	n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
	n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
	n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
	n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
	n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
	n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
	n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
	n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
	n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
	n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
	n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
	n3852, n3853, n3854, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
	n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
	n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
	n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
	n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
	n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
	n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
	n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
	n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
	n3974, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
	n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3995, n3996,
	n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4007,
	n4008, n4009, n4011, n4012, n4019, n4020, n4021, n4022, n4023, n4024,
	n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
	n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
	n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
	n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
	n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
	n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
	n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
	n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
	n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
	n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
	n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
	n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
	n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
	n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
	n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
	n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
	n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
	n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
	n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
	n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
	n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
	n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
	n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
	n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
	n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
	n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
	n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
	n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
	n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
	n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
	n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
	n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
	n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
	n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
	n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
	n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
	n4385, n4386, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
	n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
	n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
	n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
	n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
	n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
	n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
	n4456, n4457, n4458, n554, n555, n556, n557, n558, n559, n560, n561, n562,
	n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
	n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585, n586,
	n587, n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
	n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609, n610,
	n611, n612, n613, n614, n615, n616, n617, n618, n619, n620, n621, n622,
	n623, n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
	n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
	n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657, n658,
	n659, n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
	n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
	n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
	n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n707,
	n708, n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
	n720, n721, n722, n724, n725, n726, n728, n729, n731, n732, n733, n734,
	n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746,
	n747, n748, n749, n750, n752, n753, n755, n756, n757, n758, n759, n760,
	n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
	n773, n775, n776, n777, n778, n779, n780, n782, n783, n784, n785, n786,
	n787, n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
	n800, n801, n802, n803, n804, n805, n807, n808, n809, n810, n811, n812,
	n813, n815, n816, n817, n818, n820, n822, n823, n824, n825, n826, n827,
	n829, n831, n832, n833, n834, n835, n836, n837, n840, n841, n842, n843,
	n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
	n857, n859, n860, n861, n862, n863, n865, n866, n867, n868, n870, n871,
	n872, n873, n878, n879, n881, n882, n883, n884, n886, n887, n888, n889,
	n892, n895, n896, n909, n910, n911, n912, n913, n914, n915, n916, n917,
	n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
	n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940, n941,
	n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
	n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
	n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976, n977,
	n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
	n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, net148858,
	net148863, net148865, net148913, net148915, net148916, net149236, net149679,
	net149680, net149681, net150625, net150626, net150785, net151343, net151366,
	net152024, net152025, opcode_of_MEM_0, opcode_of_MEM_1, opcode_of_MEM_2,
	opcode_of_MEM_3, opcode_of_MEM_4, opcode_of_MEM_5, opcode_of_MEM_reg_0__m2s,
	opcode_of_MEM_reg_1__m2s, opcode_of_MEM_reg_2__m2s, opcode_of_MEM_reg_3__m2s,
	opcode_of_MEM_reg_4__m2s, opcode_of_MEM_reg_5__m2s, opcode_of_WB_5, opcode_of_WB_reg_0__m2s,
	opcode_of_WB_reg_1__m2s, opcode_of_WB_reg_2__m2s, opcode_of_WB_reg_3__m2s,
	opcode_of_WB_reg_4__m2s, opcode_of_WB_reg_5__m2s, rd_addr_reg_0__m2s,
	rd_addr_reg_1__m2s, rd_addr_reg_2__m2s, rd_addr_reg_3__m2s, rd_addr_reg_4__m2s,
	reg_dst_of_EX_0, reg_dst_of_EX_1, reg_dst_of_EX_2, reg_dst_of_EX_3, reg_dst_of_EX_4,
	reg_dst_of_MEM_0, reg_dst_of_MEM_1, reg_dst_of_MEM_2, reg_dst_of_MEM_3,
	reg_dst_of_MEM_4, reg_dst_of_MEM_reg_0__m2s, reg_dst_of_MEM_reg_1__m2s,
	reg_dst_of_MEM_reg_2__m2s, reg_dst_of_MEM_reg_3__m2s, reg_dst_of_MEM_reg_4__m2s,
	reg_dst_reg__m2s, reg_out_A_reg_0__m2s, reg_out_A_reg_10__m2s, reg_out_A_reg_11__m2s,
	reg_out_A_reg_12__m2s, reg_out_A_reg_13__m2s, reg_out_A_reg_14__m2s, reg_out_A_reg_15__m2s,
	reg_out_A_reg_16__m2s, reg_out_A_reg_17__m2s, reg_out_A_reg_18__m2s, reg_out_A_reg_19__m2s,
	reg_out_A_reg_1__m2s, reg_out_A_reg_20__m2s, reg_out_A_reg_21__m2s, reg_out_A_reg_22__m2s,
	reg_out_A_reg_23__m2s, reg_out_A_reg_24__m2s, reg_out_A_reg_25__m2s, reg_out_A_reg_26__m2s,
	reg_out_A_reg_27__m2s, reg_out_A_reg_28__m2s, reg_out_A_reg_29__m2s, reg_out_A_reg_2__m2s,
	reg_out_A_reg_30__m2s, reg_out_A_reg_31__m2s, reg_out_A_reg_3__m2s, reg_out_A_reg_4__m2s,
	reg_out_A_reg_5__m2s, reg_out_A_reg_6__m2s, reg_out_A_reg_7__m2s, reg_out_A_reg_8__m2s,
	reg_out_A_reg_9__m2s, reg_out_B_reg_0__m2s, reg_out_B_reg_10__m2s, reg_out_B_reg_11__m2s,
	reg_out_B_reg_12__m2s, reg_out_B_reg_13__m2s, reg_out_B_reg_14__m2s, reg_out_B_reg_15__m2s,
	reg_out_B_reg_16__m2s, reg_out_B_reg_17__m2s, reg_out_B_reg_18__m2s, reg_out_B_reg_19__m2s,
	reg_out_B_reg_1__m2s, reg_out_B_reg_20__m2s, reg_out_B_reg_21__m2s, reg_out_B_reg_22__m2s,
	reg_out_B_reg_23__m2s, reg_out_B_reg_24__m2s, reg_out_B_reg_25__m2s, reg_out_B_reg_26__m2s,
	reg_out_B_reg_27__m2s, reg_out_B_reg_28__m2s, reg_out_B_reg_29__m2s, reg_out_B_reg_2__m2s,
	reg_out_B_reg_30__m2s, reg_out_B_reg_31__m2s, reg_out_B_reg_3__m2s, reg_out_B_reg_4__m2s,
	reg_out_B_reg_5__m2s, reg_out_B_reg_6__m2s, reg_out_B_reg_7__m2s, reg_out_B_reg_8__m2s,
	reg_out_B_reg_9__m2s, reg_write_reg__m2s, rt_addr_reg_0__m2s, rt_addr_reg_1__m2s,
	rt_addr_reg_2__m2s, rt_addr_reg_3__m2s, rt_addr_reg_4__m2s, slot_num_0,
	slot_num_1, slot_num_reg_0__m2s, slot_num_reg_1__m2s, stall_reg__m2s;

	assign stall = test_so;

	DLX_sync_MUX_OP_32_5_32_2_test_1 C440 ( .D0_31(_RegFile_0__0), .D0_30(_RegFile_0__1),
		.D0_29(_RegFile_0__2), .D0_28(_RegFile_0__3), .D0_27(_RegFile_0__4),
		.D0_26(_RegFile_0__5), .D0_25(_RegFile_0__6), .D0_24(_RegFile_0__7),
		.D0_23(_RegFile_0__8), .D0_22(_RegFile_0__9), .D0_21(_RegFile_0__10),
		.D0_20(_RegFile_0__11), .D0_19(_RegFile_0__12), .D0_18(_RegFile_0__13),
		.D0_17(_RegFile_0__14), .D0_16(_RegFile_0__15), .D0_15(_RegFile_0__16),
		.D0_14(_RegFile_0__17), .D0_13(_RegFile_0__18), .D0_12(_RegFile_0__19),
		.D0_11(_RegFile_0__20), .D0_10(_RegFile_0__21), .D0_9(_RegFile_0__22),
		.D0_8(_RegFile_0__23), .D0_7(_RegFile_0__24), .D0_6(_RegFile_0__25),
		.D0_5(_RegFile_0__26), .D0_4(_RegFile_0__27), .D0_3(_RegFile_0__28),
		.D0_2(_RegFile_0__29), .D0_1(_RegFile_0__30), .D0_0(_RegFile_0__31),
		.D1_31(_RegFile_1__0), .D1_30(_RegFile_1__1), .D1_29(_RegFile_1__2),
		.D1_28(_RegFile_1__3), .D1_27(_RegFile_1__4), .D1_26(_RegFile_1__5),
		.D1_25(_RegFile_1__6), .D1_24(_RegFile_1__7), .D1_23(_RegFile_1__8),
		.D1_22(_RegFile_1__9), .D1_21(_RegFile_1__10), .D1_20(_RegFile_1__11),
		.D1_19(_RegFile_1__12), .D1_18(_RegFile_1__13), .D1_17(_RegFile_1__14),
		.D1_16(_RegFile_1__15), .D1_15(_RegFile_1__16), .D1_14(_RegFile_1__17),
		.D1_13(_RegFile_1__18), .D1_12(_RegFile_1__19), .D1_11(_RegFile_1__20),
		.D1_10(_RegFile_1__21), .D1_9(_RegFile_1__22), .D1_8(_RegFile_1__23),
		.D1_7(_RegFile_1__24), .D1_6(_RegFile_1__25), .D1_5(_RegFile_1__26),
		.D1_4(_RegFile_1__27), .D1_3(_RegFile_1__28), .D1_2(_RegFile_1__29),
		.D1_1(_RegFile_1__30), .D1_0(_RegFile_1__31), .D2_31(_RegFile_2__0),
		.D2_30(_RegFile_2__1), .D2_29(_RegFile_2__2), .D2_28(_RegFile_2__3),
		.D2_27(_RegFile_2__4), .D2_26(_RegFile_2__5), .D2_25(_RegFile_2__6),
		.D2_24(_RegFile_2__7), .D2_23(_RegFile_2__8), .D2_22(_RegFile_2__9),
		.D2_21(_RegFile_2__10), .D2_20(_RegFile_2__11), .D2_19(_RegFile_2__12),
		.D2_18(_RegFile_2__13), .D2_17(_RegFile_2__14), .D2_16(_RegFile_2__15),
		.D2_15(_RegFile_2__16), .D2_14(_RegFile_2__17), .D2_13(_RegFile_2__18),
		.D2_12(_RegFile_2__19), .D2_11(_RegFile_2__20), .D2_10(_RegFile_2__21),
		.D2_9(_RegFile_2__22), .D2_8(_RegFile_2__23), .D2_7(_RegFile_2__24),
		.D2_6(_RegFile_2__25), .D2_5(_RegFile_2__26), .D2_4(_RegFile_2__27),
		.D2_3(_RegFile_2__28), .D2_2(_RegFile_2__29), .D2_1(_RegFile_2__30),
		.D2_0(_RegFile_2__31), .D3_31(_RegFile_3__0), .D3_30(_RegFile_3__1),
		.D3_29(_RegFile_3__2), .D3_28(_RegFile_3__3), .D3_27(_RegFile_3__4),
		.D3_26(_RegFile_3__5), .D3_25(_RegFile_3__6), .D3_24(_RegFile_3__7),
		.D3_23(_RegFile_3__8), .D3_22(_RegFile_3__9), .D3_21(_RegFile_3__10),
		.D3_20(_RegFile_3__11), .D3_19(_RegFile_3__12), .D3_18(_RegFile_3__13),
		.D3_17(_RegFile_3__14), .D3_16(_RegFile_3__15), .D3_15(_RegFile_3__16),
		.D3_14(_RegFile_3__17), .D3_13(_RegFile_3__18), .D3_12(_RegFile_3__19),
		.D3_11(_RegFile_3__20), .D3_10(_RegFile_3__21), .D3_9(_RegFile_3__22),
		.D3_8(_RegFile_3__23), .D3_7(_RegFile_3__24), .D3_6(_RegFile_3__25),
		.D3_5(_RegFile_3__26), .D3_4(_RegFile_3__27), .D3_3(_RegFile_3__28),
		.D3_2(_RegFile_3__29), .D3_1(_RegFile_3__30), .D3_0(_RegFile_3__31),
		.D4_31(_RegFile_4__0), .D4_30(_RegFile_4__1), .D4_29(_RegFile_4__2),
		.D4_28(_RegFile_4__3), .D4_27(_RegFile_4__4), .D4_26(_RegFile_4__5),
		.D4_25(_RegFile_4__6), .D4_24(_RegFile_4__7), .D4_23(_RegFile_4__8),
		.D4_22(_RegFile_4__9), .D4_21(_RegFile_4__10), .D4_20(_RegFile_4__11),
		.D4_19(_RegFile_4__12), .D4_18(_RegFile_4__13), .D4_17(_RegFile_4__14),
		.D4_16(_RegFile_4__15), .D4_15(_RegFile_4__16), .D4_14(_RegFile_4__17),
		.D4_13(_RegFile_4__18), .D4_12(_RegFile_4__19), .D4_11(_RegFile_4__20),
		.D4_10(_RegFile_4__21), .D4_9(_RegFile_4__22), .D4_8(_RegFile_4__23),
		.D4_7(_RegFile_4__24), .D4_6(_RegFile_4__25), .D4_5(_RegFile_4__26),
		.D4_4(_RegFile_4__27), .D4_3(_RegFile_4__28), .D4_2(_RegFile_4__29),
		.D4_1(_RegFile_4__30), .D4_0(_RegFile_4__31), .D5_31(_RegFile_5__0),
		.D5_30(_RegFile_5__1), .D5_29(_RegFile_5__2), .D5_28(_RegFile_5__3),
		.D5_27(_RegFile_5__4), .D5_26(_RegFile_5__5), .D5_25(_RegFile_5__6),
		.D5_24(_RegFile_5__7), .D5_23(_RegFile_5__8), .D5_22(_RegFile_5__9),
		.D5_21(_RegFile_5__10), .D5_20(_RegFile_5__11), .D5_19(_RegFile_5__12),
		.D5_18(_RegFile_5__13), .D5_17(_RegFile_5__14), .D5_16(_RegFile_5__15),
		.D5_15(_RegFile_5__16), .D5_14(_RegFile_5__17), .D5_13(_RegFile_5__18),
		.D5_12(_RegFile_5__19), .D5_11(_RegFile_5__20), .D5_10(_RegFile_5__21),
		.D5_9(_RegFile_5__22), .D5_8(_RegFile_5__23), .D5_7(_RegFile_5__24),
		.D5_6(_RegFile_5__25), .D5_5(_RegFile_5__26), .D5_4(_RegFile_5__27),
		.D5_3(_RegFile_5__28), .D5_2(_RegFile_5__29), .D5_1(_RegFile_5__30),
		.D5_0(_RegFile_5__31), .D6_31(_RegFile_6__0), .D6_30(_RegFile_6__1),
		.D6_29(_RegFile_6__2), .D6_28(_RegFile_6__3), .D6_27(_RegFile_6__4),
		.D6_26(_RegFile_6__5), .D6_25(_RegFile_6__6), .D6_24(_RegFile_6__7),
		.D6_23(_RegFile_6__8), .D6_22(_RegFile_6__9), .D6_21(_RegFile_6__10),
		.D6_20(_RegFile_6__11), .D6_19(_RegFile_6__12), .D6_18(_RegFile_6__13),
		.D6_17(_RegFile_6__14), .D6_16(_RegFile_6__15), .D6_15(_RegFile_6__16),
		.D6_14(_RegFile_6__17), .D6_13(_RegFile_6__18), .D6_12(_RegFile_6__19),
		.D6_11(_RegFile_6__20), .D6_10(_RegFile_6__21), .D6_9(_RegFile_6__22),
		.D6_8(_RegFile_6__23), .D6_7(_RegFile_6__24), .D6_6(_RegFile_6__25),
		.D6_5(_RegFile_6__26), .D6_4(_RegFile_6__27), .D6_3(_RegFile_6__28),
		.D6_2(_RegFile_6__29), .D6_1(_RegFile_6__30), .D6_0(_RegFile_6__31),
		.D7_31(_RegFile_7__0), .D7_30(_RegFile_7__1), .D7_29(_RegFile_7__2),
		.D7_28(_RegFile_7__3), .D7_27(_RegFile_7__4), .D7_26(_RegFile_7__5),
		.D7_25(_RegFile_7__6), .D7_24(_RegFile_7__7), .D7_23(_RegFile_7__8),
		.D7_22(_RegFile_7__9), .D7_21(_RegFile_7__10), .D7_20(_RegFile_7__11),
		.D7_19(_RegFile_7__12), .D7_18(_RegFile_7__13), .D7_17(_RegFile_7__14),
		.D7_16(_RegFile_7__15), .D7_15(_RegFile_7__16), .D7_14(_RegFile_7__17),
		.D7_13(_RegFile_7__18), .D7_12(_RegFile_7__19), .D7_11(_RegFile_7__20),
		.D7_10(_RegFile_7__21), .D7_9(_RegFile_7__22), .D7_8(_RegFile_7__23),
		.D7_7(_RegFile_7__24), .D7_6(_RegFile_7__25), .D7_5(_RegFile_7__26),
		.D7_4(_RegFile_7__27), .D7_3(_RegFile_7__28), .D7_2(_RegFile_7__29),
		.D7_1(_RegFile_7__30), .D7_0(_RegFile_7__31), .D8_31(_RegFile_8__0),
		.D8_30(_RegFile_8__1), .D8_29(_RegFile_8__2), .D8_28(_RegFile_8__3),
		.D8_27(_RegFile_8__4), .D8_26(_RegFile_8__5), .D8_25(_RegFile_8__6),
		.D8_24(_RegFile_8__7), .D8_23(_RegFile_8__8), .D8_22(_RegFile_8__9),
		.D8_21(_RegFile_8__10), .D8_20(_RegFile_8__11), .D8_19(_RegFile_8__12),
		.D8_18(_RegFile_8__13), .D8_17(_RegFile_8__14), .D8_16(_RegFile_8__15),
		.D8_15(_RegFile_8__16), .D8_14(_RegFile_8__17), .D8_13(_RegFile_8__18),
		.D8_12(_RegFile_8__19), .D8_11(_RegFile_8__20), .D8_10(_RegFile_8__21),
		.D8_9(_RegFile_8__22), .D8_8(_RegFile_8__23), .D8_7(_RegFile_8__24),
		.D8_6(_RegFile_8__25), .D8_5(_RegFile_8__26), .D8_4(_RegFile_8__27),
		.D8_3(_RegFile_8__28), .D8_2(_RegFile_8__29), .D8_1(_RegFile_8__30),
		.D8_0(_RegFile_8__31), .D9_31(_RegFile_9__0), .D9_30(_RegFile_9__1),
		.D9_29(_RegFile_9__2), .D9_28(_RegFile_9__3), .D9_27(_RegFile_9__4),
		.D9_26(_RegFile_9__5), .D9_25(_RegFile_9__6), .D9_24(_RegFile_9__7),
		.D9_23(_RegFile_9__8), .D9_22(_RegFile_9__9), .D9_21(_RegFile_9__10),
		.D9_20(_RegFile_9__11), .D9_19(_RegFile_9__12), .D9_18(_RegFile_9__13),
		.D9_17(_RegFile_9__14), .D9_16(_RegFile_9__15), .D9_15(_RegFile_9__16),
		.D9_14(_RegFile_9__17), .D9_13(_RegFile_9__18), .D9_12(_RegFile_9__19),
		.D9_11(_RegFile_9__20), .D9_10(_RegFile_9__21), .D9_9(_RegFile_9__22),
		.D9_8(_RegFile_9__23), .D9_7(_RegFile_9__24), .D9_6(_RegFile_9__25),
		.D9_5(_RegFile_9__26), .D9_4(_RegFile_9__27), .D9_3(_RegFile_9__28),
		.D9_2(_RegFile_9__29), .D9_1(_RegFile_9__30), .D9_0(_RegFile_9__31),
		.D10_31(_RegFile_10__0), .D10_30(_RegFile_10__1), .D10_29(_RegFile_10__2),
		.D10_28(_RegFile_10__3), .D10_27(_RegFile_10__4), .D10_26(_RegFile_10__5),
		.D10_25(_RegFile_10__6), .D10_24(_RegFile_10__7), .D10_23(_RegFile_10__8),
		.D10_22(_RegFile_10__9), .D10_21(_RegFile_10__10), .D10_20(_RegFile_10__11),
		.D10_19(_RegFile_10__12), .D10_18(_RegFile_10__13), .D10_17(_RegFile_10__14),
		.D10_16(_RegFile_10__15), .D10_15(_RegFile_10__16), .D10_14(_RegFile_10__17),
		.D10_13(_RegFile_10__18), .D10_12(_RegFile_10__19), .D10_11(_RegFile_10__20),
		.D10_10(_RegFile_10__21), .D10_9(_RegFile_10__22), .D10_8(_RegFile_10__23),
		.D10_7(_RegFile_10__24), .D10_6(_RegFile_10__25), .D10_5(_RegFile_10__26),
		.D10_4(_RegFile_10__27), .D10_3(_RegFile_10__28), .D10_2(_RegFile_10__29),
		.D10_1(_RegFile_10__30), .D10_0(_RegFile_10__31), .D11_31(_RegFile_11__0),
		.D11_30(_RegFile_11__1), .D11_29(_RegFile_11__2), .D11_28(_RegFile_11__3),
		.D11_27(_RegFile_11__4), .D11_26(_RegFile_11__5), .D11_25(_RegFile_11__6),
		.D11_24(_RegFile_11__7), .D11_23(_RegFile_11__8), .D11_22(_RegFile_11__9),
		.D11_21(_RegFile_11__10), .D11_20(_RegFile_11__11), .D11_19(_RegFile_11__12),
		.D11_18(_RegFile_11__13), .D11_17(_RegFile_11__14), .D11_16(_RegFile_11__15),
		.D11_15(_RegFile_11__16), .D11_14(_RegFile_11__17), .D11_13(_RegFile_11__18),
		.D11_12(_RegFile_11__19), .D11_11(_RegFile_11__20), .D11_10(_RegFile_11__21),
		.D11_9(_RegFile_11__22), .D11_8(_RegFile_11__23), .D11_7(_RegFile_11__24),
		.D11_6(_RegFile_11__25), .D11_5(_RegFile_11__26), .D11_4(_RegFile_11__27),
		.D11_3(_RegFile_11__28), .D11_2(_RegFile_11__29), .D11_1(_RegFile_11__30),
		.D11_0(_RegFile_11__31), .D12_31(_RegFile_12__0), .D12_30(_RegFile_12__1),
		.D12_29(_RegFile_12__2), .D12_28(_RegFile_12__3), .D12_27(_RegFile_12__4),
		.D12_26(_RegFile_12__5), .D12_25(_RegFile_12__6), .D12_24(_RegFile_12__7),
		.D12_23(_RegFile_12__8), .D12_22(_RegFile_12__9), .D12_21(_RegFile_12__10),
		.D12_20(_RegFile_12__11), .D12_19(_RegFile_12__12), .D12_18(_RegFile_12__13),
		.D12_17(_RegFile_12__14), .D12_16(_RegFile_12__15), .D12_15(_RegFile_12__16),
		.D12_14(_RegFile_12__17), .D12_13(_RegFile_12__18), .D12_12(_RegFile_12__19),
		.D12_11(_RegFile_12__20), .D12_10(_RegFile_12__21), .D12_9(_RegFile_12__22),
		.D12_8(_RegFile_12__23), .D12_7(_RegFile_12__24), .D12_6(_RegFile_12__25),
		.D12_5(_RegFile_12__26), .D12_4(_RegFile_12__27), .D12_3(_RegFile_12__28),
		.D12_2(_RegFile_12__29), .D12_1(_RegFile_12__30), .D12_0(_RegFile_12__31),
		.D13_31(_RegFile_13__0), .D13_30(_RegFile_13__1), .D13_29(_RegFile_13__2),
		.D13_28(_RegFile_13__3), .D13_27(_RegFile_13__4), .D13_26(_RegFile_13__5),
		.D13_25(_RegFile_13__6), .D13_24(_RegFile_13__7), .D13_23(_RegFile_13__8),
		.D13_22(_RegFile_13__9), .D13_21(_RegFile_13__10), .D13_20(_RegFile_13__11),
		.D13_19(_RegFile_13__12), .D13_18(_RegFile_13__13), .D13_17(_RegFile_13__14),
		.D13_16(_RegFile_13__15), .D13_15(_RegFile_13__16), .D13_14(_RegFile_13__17),
		.D13_13(_RegFile_13__18), .D13_12(_RegFile_13__19), .D13_11(_RegFile_13__20),
		.D13_10(_RegFile_13__21), .D13_9(_RegFile_13__22), .D13_8(_RegFile_13__23),
		.D13_7(_RegFile_13__24), .D13_6(_RegFile_13__25), .D13_5(_RegFile_13__26),
		.D13_4(_RegFile_13__27), .D13_3(_RegFile_13__28), .D13_2(_RegFile_13__29),
		.D13_1(_RegFile_13__30), .D13_0(_RegFile_13__31), .D14_31(_RegFile_14__0),
		.D14_30(_RegFile_14__1), .D14_29(_RegFile_14__2), .D14_28(_RegFile_14__3),
		.D14_27(_RegFile_14__4), .D14_26(_RegFile_14__5), .D14_25(_RegFile_14__6),
		.D14_24(_RegFile_14__7), .D14_23(_RegFile_14__8), .D14_22(_RegFile_14__9),
		.D14_21(_RegFile_14__10), .D14_20(_RegFile_14__11), .D14_19(_RegFile_14__12),
		.D14_18(_RegFile_14__13), .D14_17(_RegFile_14__14), .D14_16(_RegFile_14__15),
		.D14_15(_RegFile_14__16), .D14_14(_RegFile_14__17), .D14_13(_RegFile_14__18),
		.D14_12(_RegFile_14__19), .D14_11(_RegFile_14__20), .D14_10(_RegFile_14__21),
		.D14_9(_RegFile_14__22), .D14_8(_RegFile_14__23), .D14_7(_RegFile_14__24),
		.D14_6(_RegFile_14__25), .D14_5(_RegFile_14__26), .D14_4(_RegFile_14__27),
		.D14_3(_RegFile_14__28), .D14_2(_RegFile_14__29), .D14_1(_RegFile_14__30),
		.D14_0(_RegFile_14__31), .D15_31(_RegFile_15__0), .D15_30(_RegFile_15__1),
		.D15_29(_RegFile_15__2), .D15_28(_RegFile_15__3), .D15_27(_RegFile_15__4),
		.D15_26(_RegFile_15__5), .D15_25(_RegFile_15__6), .D15_24(_RegFile_15__7),
		.D15_23(_RegFile_15__8), .D15_22(_RegFile_15__9), .D15_21(_RegFile_15__10),
		.D15_20(_RegFile_15__11), .D15_19(_RegFile_15__12), .D15_18(_RegFile_15__13),
		.D15_17(_RegFile_15__14), .D15_16(_RegFile_15__15), .D15_15(_RegFile_15__16),
		.D15_14(_RegFile_15__17), .D15_13(_RegFile_15__18), .D15_12(_RegFile_15__19),
		.D15_11(_RegFile_15__20), .D15_10(_RegFile_15__21), .D15_9(_RegFile_15__22),
		.D15_8(_RegFile_15__23), .D15_7(_RegFile_15__24), .D15_6(_RegFile_15__25),
		.D15_5(_RegFile_15__26), .D15_4(_RegFile_15__27), .D15_3(_RegFile_15__28),
		.D15_2(_RegFile_15__29), .D15_1(_RegFile_15__30), .D15_0(_RegFile_15__31),
		.D16_31(_RegFile_16__0), .D16_30(_RegFile_16__1), .D16_29(_RegFile_16__2),
		.D16_28(_RegFile_16__3), .D16_27(_RegFile_16__4), .D16_26(_RegFile_16__5),
		.D16_25(_RegFile_16__6), .D16_24(_RegFile_16__7), .D16_23(_RegFile_16__8),
		.D16_22(_RegFile_16__9), .D16_21(_RegFile_16__10), .D16_20(_RegFile_16__11),
		.D16_19(_RegFile_16__12), .D16_18(_RegFile_16__13), .D16_17(_RegFile_16__14),
		.D16_16(_RegFile_16__15), .D16_15(_RegFile_16__16), .D16_14(_RegFile_16__17),
		.D16_13(_RegFile_16__18), .D16_12(_RegFile_16__19), .D16_11(_RegFile_16__20),
		.D16_10(_RegFile_16__21), .D16_9(_RegFile_16__22), .D16_8(_RegFile_16__23),
		.D16_7(_RegFile_16__24), .D16_6(_RegFile_16__25), .D16_5(_RegFile_16__26),
		.D16_4(_RegFile_16__27), .D16_3(_RegFile_16__28), .D16_2(_RegFile_16__29),
		.D16_1(_RegFile_16__30), .D16_0(_RegFile_16__31), .D17_31(_RegFile_17__0),
		.D17_30(_RegFile_17__1), .D17_29(_RegFile_17__2), .D17_28(_RegFile_17__3),
		.D17_27(_RegFile_17__4), .D17_26(_RegFile_17__5), .D17_25(_RegFile_17__6),
		.D17_24(_RegFile_17__7), .D17_23(_RegFile_17__8), .D17_22(_RegFile_17__9),
		.D17_21(_RegFile_17__10), .D17_20(_RegFile_17__11), .D17_19(_RegFile_17__12),
		.D17_18(_RegFile_17__13), .D17_17(_RegFile_17__14), .D17_16(_RegFile_17__15),
		.D17_15(_RegFile_17__16), .D17_14(_RegFile_17__17), .D17_13(_RegFile_17__18),
		.D17_12(_RegFile_17__19), .D17_11(_RegFile_17__20), .D17_10(_RegFile_17__21),
		.D17_9(_RegFile_17__22), .D17_8(_RegFile_17__23), .D17_7(_RegFile_17__24),
		.D17_6(_RegFile_17__25), .D17_5(_RegFile_17__26), .D17_4(_RegFile_17__27),
		.D17_3(_RegFile_17__28), .D17_2(_RegFile_17__29), .D17_1(_RegFile_17__30),
		.D17_0(_RegFile_17__31), .D18_31(_RegFile_18__0), .D18_30(_RegFile_18__1),
		.D18_29(_RegFile_18__2), .D18_28(_RegFile_18__3), .D18_27(_RegFile_18__4),
		.D18_26(_RegFile_18__5), .D18_25(_RegFile_18__6), .D18_24(_RegFile_18__7),
		.D18_23(_RegFile_18__8), .D18_22(_RegFile_18__9), .D18_21(_RegFile_18__10),
		.D18_20(_RegFile_18__11), .D18_19(_RegFile_18__12), .D18_18(_RegFile_18__13),
		.D18_17(_RegFile_18__14), .D18_16(_RegFile_18__15), .D18_15(_RegFile_18__16),
		.D18_14(_RegFile_18__17), .D18_13(_RegFile_18__18), .D18_12(_RegFile_18__19),
		.D18_11(_RegFile_18__20), .D18_10(_RegFile_18__21), .D18_9(_RegFile_18__22),
		.D18_8(_RegFile_18__23), .D18_7(_RegFile_18__24), .D18_6(_RegFile_18__25),
		.D18_5(_RegFile_18__26), .D18_4(_RegFile_18__27), .D18_3(_RegFile_18__28),
		.D18_2(_RegFile_18__29), .D18_1(_RegFile_18__30), .D18_0(_RegFile_18__31),
		.D19_31(_RegFile_19__0), .D19_30(_RegFile_19__1), .D19_29(_RegFile_19__2),
		.D19_28(_RegFile_19__3), .D19_27(_RegFile_19__4), .D19_26(_RegFile_19__5),
		.D19_25(_RegFile_19__6), .D19_24(_RegFile_19__7), .D19_23(_RegFile_19__8),
		.D19_22(_RegFile_19__9), .D19_21(_RegFile_19__10), .D19_20(_RegFile_19__11),
		.D19_19(_RegFile_19__12), .D19_18(_RegFile_19__13), .D19_17(_RegFile_19__14),
		.D19_16(_RegFile_19__15), .D19_15(_RegFile_19__16), .D19_14(_RegFile_19__17),
		.D19_13(_RegFile_19__18), .D19_12(_RegFile_19__19), .D19_11(_RegFile_19__20),
		.D19_10(_RegFile_19__21), .D19_9(_RegFile_19__22), .D19_8(_RegFile_19__23),
		.D19_7(_RegFile_19__24), .D19_6(_RegFile_19__25), .D19_5(_RegFile_19__26),
		.D19_4(_RegFile_19__27), .D19_3(_RegFile_19__28), .D19_2(_RegFile_19__29),
		.D19_1(_RegFile_19__30), .D19_0(_RegFile_19__31), .D20_31(_RegFile_20__0),
		.D20_30(_RegFile_20__1), .D20_29(_RegFile_20__2), .D20_28(_RegFile_20__3),
		.D20_27(_RegFile_20__4), .D20_26(_RegFile_20__5), .D20_25(_RegFile_20__6),
		.D20_24(_RegFile_20__7), .D20_23(_RegFile_20__8), .D20_22(_RegFile_20__9),
		.D20_21(_RegFile_20__10), .D20_20(_RegFile_20__11), .D20_19(_RegFile_20__12),
		.D20_18(_RegFile_20__13), .D20_17(_RegFile_20__14), .D20_16(_RegFile_20__15),
		.D20_15(_RegFile_20__16), .D20_14(_RegFile_20__17), .D20_13(_RegFile_20__18),
		.D20_12(_RegFile_20__19), .D20_11(_RegFile_20__20), .D20_10(_RegFile_20__21),
		.D20_9(_RegFile_20__22), .D20_8(_RegFile_20__23), .D20_7(_RegFile_20__24),
		.D20_6(_RegFile_20__25), .D20_5(_RegFile_20__26), .D20_4(_RegFile_20__27),
		.D20_3(_RegFile_20__28), .D20_2(_RegFile_20__29), .D20_1(_RegFile_20__30),
		.D20_0(_RegFile_20__31), .D21_31(_RegFile_21__0), .D21_30(_RegFile_21__1),
		.D21_29(_RegFile_21__2), .D21_28(_RegFile_21__3), .D21_27(_RegFile_21__4),
		.D21_26(_RegFile_21__5), .D21_25(_RegFile_21__6), .D21_24(_RegFile_21__7),
		.D21_23(_RegFile_21__8), .D21_22(_RegFile_21__9), .D21_21(_RegFile_21__10),
		.D21_20(_RegFile_21__11), .D21_19(_RegFile_21__12), .D21_18(_RegFile_21__13),
		.D21_17(_RegFile_21__14), .D21_16(_RegFile_21__15), .D21_15(_RegFile_21__16),
		.D21_14(_RegFile_21__17), .D21_13(_RegFile_21__18), .D21_12(_RegFile_21__19),
		.D21_11(_RegFile_21__20), .D21_10(_RegFile_21__21), .D21_9(_RegFile_21__22),
		.D21_8(_RegFile_21__23), .D21_7(_RegFile_21__24), .D21_6(_RegFile_21__25),
		.D21_5(_RegFile_21__26), .D21_4(_RegFile_21__27), .D21_3(_RegFile_21__28),
		.D21_2(_RegFile_21__29), .D21_1(_RegFile_21__30), .D21_0(_RegFile_21__31),
		.D22_31(_RegFile_22__0), .D22_30(_RegFile_22__1), .D22_29(_RegFile_22__2),
		.D22_28(_RegFile_22__3), .D22_27(_RegFile_22__4), .D22_26(_RegFile_22__5),
		.D22_25(_RegFile_22__6), .D22_24(_RegFile_22__7), .D22_23(_RegFile_22__8),
		.D22_22(_RegFile_22__9), .D22_21(_RegFile_22__10), .D22_20(_RegFile_22__11),
		.D22_19(_RegFile_22__12), .D22_18(_RegFile_22__13), .D22_17(_RegFile_22__14),
		.D22_16(_RegFile_22__15), .D22_15(_RegFile_22__16), .D22_14(_RegFile_22__17),
		.D22_13(_RegFile_22__18), .D22_12(_RegFile_22__19), .D22_11(_RegFile_22__20),
		.D22_10(_RegFile_22__21), .D22_9(_RegFile_22__22), .D22_8(_RegFile_22__23),
		.D22_7(_RegFile_22__24), .D22_6(_RegFile_22__25), .D22_5(_RegFile_22__26),
		.D22_4(_RegFile_22__27), .D22_3(_RegFile_22__28), .D22_2(_RegFile_22__29),
		.D22_1(_RegFile_22__30), .D22_0(_RegFile_22__31), .D23_31(_RegFile_23__0),
		.D23_30(_RegFile_23__1), .D23_29(_RegFile_23__2), .D23_28(_RegFile_23__3),
		.D23_27(_RegFile_23__4), .D23_26(_RegFile_23__5), .D23_25(_RegFile_23__6),
		.D23_24(_RegFile_23__7), .D23_23(_RegFile_23__8), .D23_22(_RegFile_23__9),
		.D23_21(_RegFile_23__10), .D23_20(_RegFile_23__11), .D23_19(_RegFile_23__12),
		.D23_18(_RegFile_23__13), .D23_17(_RegFile_23__14), .D23_16(_RegFile_23__15),
		.D23_15(_RegFile_23__16), .D23_14(_RegFile_23__17), .D23_13(_RegFile_23__18),
		.D23_12(_RegFile_23__19), .D23_11(_RegFile_23__20), .D23_10(_RegFile_23__21),
		.D23_9(_RegFile_23__22), .D23_8(_RegFile_23__23), .D23_7(_RegFile_23__24),
		.D23_6(_RegFile_23__25), .D23_5(_RegFile_23__26), .D23_4(_RegFile_23__27),
		.D23_3(_RegFile_23__28), .D23_2(_RegFile_23__29), .D23_1(_RegFile_23__30),
		.D23_0(_RegFile_23__31), .D24_31(_RegFile_24__0), .D24_30(_RegFile_24__1),
		.D24_29(_RegFile_24__2), .D24_28(_RegFile_24__3), .D24_27(_RegFile_24__4),
		.D24_26(_RegFile_24__5), .D24_25(_RegFile_24__6), .D24_24(_RegFile_24__7),
		.D24_23(_RegFile_24__8), .D24_22(_RegFile_24__9), .D24_21(_RegFile_24__10),
		.D24_20(_RegFile_24__11), .D24_19(_RegFile_24__12), .D24_18(_RegFile_24__13),
		.D24_17(_RegFile_24__14), .D24_16(_RegFile_24__15), .D24_15(_RegFile_24__16),
		.D24_14(_RegFile_24__17), .D24_13(_RegFile_24__18), .D24_12(_RegFile_24__19),
		.D24_11(_RegFile_24__20), .D24_10(_RegFile_24__21), .D24_9(_RegFile_24__22),
		.D24_8(_RegFile_24__23), .D24_7(_RegFile_24__24), .D24_6(_RegFile_24__25),
		.D24_5(_RegFile_24__26), .D24_4(_RegFile_24__27), .D24_3(_RegFile_24__28),
		.D24_2(_RegFile_24__29), .D24_1(_RegFile_24__30), .D24_0(_RegFile_24__31),
		.D25_31(_RegFile_25__0), .D25_30(_RegFile_25__1), .D25_29(_RegFile_25__2),
		.D25_28(_RegFile_25__3), .D25_27(_RegFile_25__4), .D25_26(_RegFile_25__5),
		.D25_25(_RegFile_25__6), .D25_24(_RegFile_25__7), .D25_23(_RegFile_25__8),
		.D25_22(_RegFile_25__9), .D25_21(_RegFile_25__10), .D25_20(_RegFile_25__11),
		.D25_19(_RegFile_25__12), .D25_18(_RegFile_25__13), .D25_17(_RegFile_25__14),
		.D25_16(_RegFile_25__15), .D25_15(_RegFile_25__16), .D25_14(_RegFile_25__17),
		.D25_13(_RegFile_25__18), .D25_12(_RegFile_25__19), .D25_11(_RegFile_25__20),
		.D25_10(_RegFile_25__21), .D25_9(_RegFile_25__22), .D25_8(_RegFile_25__23),
		.D25_7(_RegFile_25__24), .D25_6(_RegFile_25__25), .D25_5(_RegFile_25__26),
		.D25_4(_RegFile_25__27), .D25_3(_RegFile_25__28), .D25_2(_RegFile_25__29),
		.D25_1(_RegFile_25__30), .D25_0(_RegFile_25__31), .D26_31(_RegFile_26__0),
		.D26_30(_RegFile_26__1), .D26_29(_RegFile_26__2), .D26_28(_RegFile_26__3),
		.D26_27(_RegFile_26__4), .D26_26(_RegFile_26__5), .D26_25(_RegFile_26__6),
		.D26_24(_RegFile_26__7), .D26_23(_RegFile_26__8), .D26_22(_RegFile_26__9),
		.D26_21(_RegFile_26__10), .D26_20(_RegFile_26__11), .D26_19(_RegFile_26__12),
		.D26_18(_RegFile_26__13), .D26_17(_RegFile_26__14), .D26_16(_RegFile_26__15),
		.D26_15(_RegFile_26__16), .D26_14(_RegFile_26__17), .D26_13(_RegFile_26__18),
		.D26_12(_RegFile_26__19), .D26_11(_RegFile_26__20), .D26_10(_RegFile_26__21),
		.D26_9(_RegFile_26__22), .D26_8(_RegFile_26__23), .D26_7(_RegFile_26__24),
		.D26_6(_RegFile_26__25), .D26_5(_RegFile_26__26), .D26_4(_RegFile_26__27),
		.D26_3(_RegFile_26__28), .D26_2(_RegFile_26__29), .D26_1(_RegFile_26__30),
		.D26_0(_RegFile_26__31), .D27_31(_RegFile_27__0), .D27_30(_RegFile_27__1),
		.D27_29(_RegFile_27__2), .D27_28(_RegFile_27__3), .D27_27(_RegFile_27__4),
		.D27_26(_RegFile_27__5), .D27_25(_RegFile_27__6), .D27_24(_RegFile_27__7),
		.D27_23(_RegFile_27__8), .D27_22(_RegFile_27__9), .D27_21(_RegFile_27__10),
		.D27_20(_RegFile_27__11), .D27_19(_RegFile_27__12), .D27_18(_RegFile_27__13),
		.D27_17(_RegFile_27__14), .D27_16(_RegFile_27__15), .D27_15(_RegFile_27__16),
		.D27_14(_RegFile_27__17), .D27_13(_RegFile_27__18), .D27_12(_RegFile_27__19),
		.D27_11(_RegFile_27__20), .D27_10(_RegFile_27__21), .D27_9(_RegFile_27__22),
		.D27_8(_RegFile_27__23), .D27_7(_RegFile_27__24), .D27_6(_RegFile_27__25),
		.D27_5(_RegFile_27__26), .D27_4(_RegFile_27__27), .D27_3(_RegFile_27__28),
		.D27_2(_RegFile_27__29), .D27_1(_RegFile_27__30), .D27_0(_RegFile_27__31),
		.D28_31(_RegFile_28__0), .D28_30(_RegFile_28__1), .D28_29(_RegFile_28__2),
		.D28_28(_RegFile_28__3), .D28_27(_RegFile_28__4), .D28_26(_RegFile_28__5),
		.D28_25(_RegFile_28__6), .D28_24(_RegFile_28__7), .D28_23(_RegFile_28__8),
		.D28_22(_RegFile_28__9), .D28_21(_RegFile_28__10), .D28_20(_RegFile_28__11),
		.D28_19(_RegFile_28__12), .D28_18(_RegFile_28__13), .D28_17(_RegFile_28__14),
		.D28_16(_RegFile_28__15), .D28_15(_RegFile_28__16), .D28_14(_RegFile_28__17),
		.D28_13(_RegFile_28__18), .D28_12(_RegFile_28__19), .D28_11(_RegFile_28__20),
		.D28_10(_RegFile_28__21), .D28_9(_RegFile_28__22), .D28_8(_RegFile_28__23),
		.D28_7(_RegFile_28__24), .D28_6(_RegFile_28__25), .D28_5(_RegFile_28__26),
		.D28_4(_RegFile_28__27), .D28_3(_RegFile_28__28), .D28_2(_RegFile_28__29),
		.D28_1(_RegFile_28__30), .D28_0(_RegFile_28__31), .D29_31(_RegFile_29__0),
		.D29_30(_RegFile_29__1), .D29_29(_RegFile_29__2), .D29_28(_RegFile_29__3),
		.D29_27(_RegFile_29__4), .D29_26(_RegFile_29__5), .D29_25(_RegFile_29__6),
		.D29_24(_RegFile_29__7), .D29_23(_RegFile_29__8), .D29_22(_RegFile_29__9),
		.D29_21(_RegFile_29__10), .D29_20(_RegFile_29__11), .D29_19(_RegFile_29__12),
		.D29_18(_RegFile_29__13), .D29_17(_RegFile_29__14), .D29_16(_RegFile_29__15),
		.D29_15(_RegFile_29__16), .D29_14(_RegFile_29__17), .D29_13(_RegFile_29__18),
		.D29_12(_RegFile_29__19), .D29_11(_RegFile_29__20), .D29_10(_RegFile_29__21),
		.D29_9(_RegFile_29__22), .D29_8(_RegFile_29__23), .D29_7(_RegFile_29__24),
		.D29_6(_RegFile_29__25), .D29_5(_RegFile_29__26), .D29_4(_RegFile_29__27),
		.D29_3(_RegFile_29__28), .D29_2(_RegFile_29__29), .D29_1(_RegFile_29__30),
		.D29_0(_RegFile_29__31), .D30_31(_RegFile_30__0), .D30_30(_RegFile_30__1),
		.D30_29(_RegFile_30__2), .D30_28(_RegFile_30__3), .D30_27(_RegFile_30__4),
		.D30_26(_RegFile_30__5), .D30_25(_RegFile_30__6), .D30_24(_RegFile_30__7),
		.D30_23(_RegFile_30__8), .D30_22(_RegFile_30__9), .D30_21(_RegFile_30__10),
		.D30_20(_RegFile_30__11), .D30_19(_RegFile_30__12), .D30_18(_RegFile_30__13),
		.D30_17(_RegFile_30__14), .D30_16(_RegFile_30__15), .D30_15(_RegFile_30__16),
		.D30_14(_RegFile_30__17), .D30_13(_RegFile_30__18), .D30_12(_RegFile_30__19),
		.D30_11(_RegFile_30__20), .D30_10(_RegFile_30__21), .D30_9(_RegFile_30__22),
		.D30_8(_RegFile_30__23), .D30_7(_RegFile_30__24), .D30_6(_RegFile_30__25),
		.D30_5(_RegFile_30__26), .D30_4(_RegFile_30__27), .D30_3(_RegFile_30__28),
		.D30_2(_RegFile_30__29), .D30_1(_RegFile_30__30), .D30_0(_RegFile_30__31),
		.D31_31(_RegFile_31__0), .D31_30(_RegFile_31__1), .D31_29(_RegFile_31__2),
		.D31_28(_RegFile_31__3), .D31_27(_RegFile_31__4), .D31_26(_RegFile_31__5),
		.D31_25(_RegFile_31__6), .D31_24(_RegFile_31__7), .D31_23(_RegFile_31__8),
		.D31_22(_RegFile_31__9), .D31_21(_RegFile_31__10), .D31_20(_RegFile_31__11),
		.D31_19(_RegFile_31__12), .D31_18(_RegFile_31__13), .D31_17(_RegFile_31__14),
		.D31_16(_RegFile_31__15), .D31_15(_RegFile_31__16), .D31_14(_RegFile_31__17),
		.D31_13(_RegFile_31__18), .D31_12(_RegFile_31__19), .D31_11(_RegFile_31__20),
		.D31_10(_RegFile_31__21), .D31_9(_RegFile_31__22), .D31_8(_RegFile_31__23),
		.D31_7(_RegFile_31__24), .D31_6(_RegFile_31__25), .D31_5(_RegFile_31__26),
		.D31_4(_RegFile_31__27), .D31_3(_RegFile_31__28), .D31_2(_RegFile_31__29),
		.D31_1(_RegFile_31__30), .D31_0(_RegFile_31__31), .S0(n804), .S1(n896),
		.S2(n694), .S3(n332), .S4(n331), .Z_31(N468), .Z_30(N467), .Z_29(N466),
		.Z_28(N465), .Z_27(N464), .Z_26(N463), .Z_25(N462), .Z_24(N461), .Z_23(N460),
		.Z_22(N459), .Z_21(N458), .Z_20(N457), .Z_19(N456), .Z_18(N455), .Z_17(N454),
		.Z_16(N453), .Z_15(N452), .Z_14(N451), .Z_13(N450), .Z_12(N449), .Z_11(N448),
		.Z_10(N447), .Z_9(N446), .Z_8(N445), .Z_7(N444), .Z_6(N443), .Z_5(N442),
		.Z_4(N441), .Z_3(N440), .Z_2(N439), .Z_1(N438), .Z_0(N437) );
	DLX_sync_MUX_OP_32_5_32_test_1 C476 ( .D0_31(_RegFile_0__0), .D0_30(_RegFile_0__1),
		.D0_29(_RegFile_0__2), .D0_28(_RegFile_0__3), .D0_27(_RegFile_0__4),
		.D0_26(_RegFile_0__5), .D0_25(_RegFile_0__6), .D0_24(_RegFile_0__7),
		.D0_23(_RegFile_0__8), .D0_22(_RegFile_0__9), .D0_21(_RegFile_0__10),
		.D0_20(_RegFile_0__11), .D0_19(_RegFile_0__12), .D0_18(_RegFile_0__13),
		.D0_17(_RegFile_0__14), .D0_16(_RegFile_0__15), .D0_15(_RegFile_0__16),
		.D0_14(_RegFile_0__17), .D0_13(_RegFile_0__18), .D0_12(_RegFile_0__19),
		.D0_11(_RegFile_0__20), .D0_10(_RegFile_0__21), .D0_9(_RegFile_0__22),
		.D0_8(_RegFile_0__23), .D0_7(_RegFile_0__24), .D0_6(_RegFile_0__25),
		.D0_5(_RegFile_0__26), .D0_4(_RegFile_0__27), .D0_3(_RegFile_0__28),
		.D0_2(_RegFile_0__29), .D0_1(_RegFile_0__30), .D0_0(_RegFile_0__31),
		.D1_31(_RegFile_1__0), .D1_30(_RegFile_1__1), .D1_29(_RegFile_1__2),
		.D1_28(_RegFile_1__3), .D1_27(_RegFile_1__4), .D1_26(_RegFile_1__5),
		.D1_25(_RegFile_1__6), .D1_24(_RegFile_1__7), .D1_23(_RegFile_1__8),
		.D1_22(_RegFile_1__9), .D1_21(_RegFile_1__10), .D1_20(_RegFile_1__11),
		.D1_19(_RegFile_1__12), .D1_18(_RegFile_1__13), .D1_17(_RegFile_1__14),
		.D1_16(_RegFile_1__15), .D1_15(_RegFile_1__16), .D1_14(_RegFile_1__17),
		.D1_13(_RegFile_1__18), .D1_12(_RegFile_1__19), .D1_11(_RegFile_1__20),
		.D1_10(_RegFile_1__21), .D1_9(_RegFile_1__22), .D1_8(_RegFile_1__23),
		.D1_7(_RegFile_1__24), .D1_6(_RegFile_1__25), .D1_5(_RegFile_1__26),
		.D1_4(_RegFile_1__27), .D1_3(_RegFile_1__28), .D1_2(_RegFile_1__29),
		.D1_1(_RegFile_1__30), .D1_0(_RegFile_1__31), .D2_31(_RegFile_2__0),
		.D2_30(_RegFile_2__1), .D2_29(_RegFile_2__2), .D2_28(_RegFile_2__3),
		.D2_27(_RegFile_2__4), .D2_26(_RegFile_2__5), .D2_25(_RegFile_2__6),
		.D2_24(_RegFile_2__7), .D2_23(_RegFile_2__8), .D2_22(_RegFile_2__9),
		.D2_21(_RegFile_2__10), .D2_20(_RegFile_2__11), .D2_19(_RegFile_2__12),
		.D2_18(_RegFile_2__13), .D2_17(_RegFile_2__14), .D2_16(_RegFile_2__15),
		.D2_15(_RegFile_2__16), .D2_14(_RegFile_2__17), .D2_13(_RegFile_2__18),
		.D2_12(_RegFile_2__19), .D2_11(_RegFile_2__20), .D2_10(_RegFile_2__21),
		.D2_9(_RegFile_2__22), .D2_8(_RegFile_2__23), .D2_7(_RegFile_2__24),
		.D2_6(_RegFile_2__25), .D2_5(_RegFile_2__26), .D2_4(_RegFile_2__27),
		.D2_3(_RegFile_2__28), .D2_2(_RegFile_2__29), .D2_1(_RegFile_2__30),
		.D2_0(_RegFile_2__31), .D3_31(_RegFile_3__0), .D3_30(_RegFile_3__1),
		.D3_29(_RegFile_3__2), .D3_28(_RegFile_3__3), .D3_27(_RegFile_3__4),
		.D3_26(_RegFile_3__5), .D3_25(_RegFile_3__6), .D3_24(_RegFile_3__7),
		.D3_23(_RegFile_3__8), .D3_22(_RegFile_3__9), .D3_21(_RegFile_3__10),
		.D3_20(_RegFile_3__11), .D3_19(_RegFile_3__12), .D3_18(_RegFile_3__13),
		.D3_17(_RegFile_3__14), .D3_16(_RegFile_3__15), .D3_15(_RegFile_3__16),
		.D3_14(_RegFile_3__17), .D3_13(_RegFile_3__18), .D3_12(_RegFile_3__19),
		.D3_11(_RegFile_3__20), .D3_10(_RegFile_3__21), .D3_9(_RegFile_3__22),
		.D3_8(_RegFile_3__23), .D3_7(_RegFile_3__24), .D3_6(_RegFile_3__25),
		.D3_5(_RegFile_3__26), .D3_4(_RegFile_3__27), .D3_3(_RegFile_3__28),
		.D3_2(_RegFile_3__29), .D3_1(_RegFile_3__30), .D3_0(_RegFile_3__31),
		.D4_31(_RegFile_4__0), .D4_30(_RegFile_4__1), .D4_29(_RegFile_4__2),
		.D4_28(_RegFile_4__3), .D4_27(_RegFile_4__4), .D4_26(_RegFile_4__5),
		.D4_25(_RegFile_4__6), .D4_24(_RegFile_4__7), .D4_23(_RegFile_4__8),
		.D4_22(_RegFile_4__9), .D4_21(_RegFile_4__10), .D4_20(_RegFile_4__11),
		.D4_19(_RegFile_4__12), .D4_18(_RegFile_4__13), .D4_17(_RegFile_4__14),
		.D4_16(_RegFile_4__15), .D4_15(_RegFile_4__16), .D4_14(_RegFile_4__17),
		.D4_13(_RegFile_4__18), .D4_12(_RegFile_4__19), .D4_11(_RegFile_4__20),
		.D4_10(_RegFile_4__21), .D4_9(_RegFile_4__22), .D4_8(_RegFile_4__23),
		.D4_7(_RegFile_4__24), .D4_6(_RegFile_4__25), .D4_5(_RegFile_4__26),
		.D4_4(_RegFile_4__27), .D4_3(_RegFile_4__28), .D4_2(_RegFile_4__29),
		.D4_1(_RegFile_4__30), .D4_0(_RegFile_4__31), .D5_31(_RegFile_5__0),
		.D5_30(_RegFile_5__1), .D5_29(_RegFile_5__2), .D5_28(_RegFile_5__3),
		.D5_27(_RegFile_5__4), .D5_26(_RegFile_5__5), .D5_25(_RegFile_5__6),
		.D5_24(_RegFile_5__7), .D5_23(_RegFile_5__8), .D5_22(_RegFile_5__9),
		.D5_21(_RegFile_5__10), .D5_20(_RegFile_5__11), .D5_19(_RegFile_5__12),
		.D5_18(_RegFile_5__13), .D5_17(_RegFile_5__14), .D5_16(_RegFile_5__15),
		.D5_15(_RegFile_5__16), .D5_14(_RegFile_5__17), .D5_13(_RegFile_5__18),
		.D5_12(_RegFile_5__19), .D5_11(_RegFile_5__20), .D5_10(_RegFile_5__21),
		.D5_9(_RegFile_5__22), .D5_8(_RegFile_5__23), .D5_7(_RegFile_5__24),
		.D5_6(_RegFile_5__25), .D5_5(_RegFile_5__26), .D5_4(_RegFile_5__27),
		.D5_3(_RegFile_5__28), .D5_2(_RegFile_5__29), .D5_1(_RegFile_5__30),
		.D5_0(_RegFile_5__31), .D6_31(_RegFile_6__0), .D6_30(_RegFile_6__1),
		.D6_29(_RegFile_6__2), .D6_28(_RegFile_6__3), .D6_27(_RegFile_6__4),
		.D6_26(_RegFile_6__5), .D6_25(_RegFile_6__6), .D6_24(_RegFile_6__7),
		.D6_23(_RegFile_6__8), .D6_22(_RegFile_6__9), .D6_21(_RegFile_6__10),
		.D6_20(_RegFile_6__11), .D6_19(_RegFile_6__12), .D6_18(_RegFile_6__13),
		.D6_17(_RegFile_6__14), .D6_16(_RegFile_6__15), .D6_15(_RegFile_6__16),
		.D6_14(_RegFile_6__17), .D6_13(_RegFile_6__18), .D6_12(_RegFile_6__19),
		.D6_11(_RegFile_6__20), .D6_10(_RegFile_6__21), .D6_9(_RegFile_6__22),
		.D6_8(_RegFile_6__23), .D6_7(_RegFile_6__24), .D6_6(_RegFile_6__25),
		.D6_5(_RegFile_6__26), .D6_4(_RegFile_6__27), .D6_3(_RegFile_6__28),
		.D6_2(_RegFile_6__29), .D6_1(_RegFile_6__30), .D6_0(_RegFile_6__31),
		.D7_31(_RegFile_7__0), .D7_30(_RegFile_7__1), .D7_29(_RegFile_7__2),
		.D7_28(_RegFile_7__3), .D7_27(_RegFile_7__4), .D7_26(_RegFile_7__5),
		.D7_25(_RegFile_7__6), .D7_24(_RegFile_7__7), .D7_23(_RegFile_7__8),
		.D7_22(_RegFile_7__9), .D7_21(_RegFile_7__10), .D7_20(_RegFile_7__11),
		.D7_19(_RegFile_7__12), .D7_18(_RegFile_7__13), .D7_17(_RegFile_7__14),
		.D7_16(_RegFile_7__15), .D7_15(_RegFile_7__16), .D7_14(_RegFile_7__17),
		.D7_13(_RegFile_7__18), .D7_12(_RegFile_7__19), .D7_11(_RegFile_7__20),
		.D7_10(_RegFile_7__21), .D7_9(_RegFile_7__22), .D7_8(_RegFile_7__23),
		.D7_7(_RegFile_7__24), .D7_6(_RegFile_7__25), .D7_5(_RegFile_7__26),
		.D7_4(_RegFile_7__27), .D7_3(_RegFile_7__28), .D7_2(_RegFile_7__29),
		.D7_1(_RegFile_7__30), .D7_0(_RegFile_7__31), .D8_31(_RegFile_8__0),
		.D8_30(_RegFile_8__1), .D8_29(_RegFile_8__2), .D8_28(_RegFile_8__3),
		.D8_27(_RegFile_8__4), .D8_26(_RegFile_8__5), .D8_25(_RegFile_8__6),
		.D8_24(_RegFile_8__7), .D8_23(_RegFile_8__8), .D8_22(_RegFile_8__9),
		.D8_21(_RegFile_8__10), .D8_20(_RegFile_8__11), .D8_19(_RegFile_8__12),
		.D8_18(_RegFile_8__13), .D8_17(_RegFile_8__14), .D8_16(_RegFile_8__15),
		.D8_15(_RegFile_8__16), .D8_14(_RegFile_8__17), .D8_13(_RegFile_8__18),
		.D8_12(_RegFile_8__19), .D8_11(_RegFile_8__20), .D8_10(_RegFile_8__21),
		.D8_9(_RegFile_8__22), .D8_8(_RegFile_8__23), .D8_7(_RegFile_8__24),
		.D8_6(_RegFile_8__25), .D8_5(_RegFile_8__26), .D8_4(_RegFile_8__27),
		.D8_3(_RegFile_8__28), .D8_2(_RegFile_8__29), .D8_1(_RegFile_8__30),
		.D8_0(_RegFile_8__31), .D9_31(_RegFile_9__0), .D9_30(_RegFile_9__1),
		.D9_29(_RegFile_9__2), .D9_28(_RegFile_9__3), .D9_27(_RegFile_9__4),
		.D9_26(_RegFile_9__5), .D9_25(_RegFile_9__6), .D9_24(_RegFile_9__7),
		.D9_23(_RegFile_9__8), .D9_22(_RegFile_9__9), .D9_21(_RegFile_9__10),
		.D9_20(_RegFile_9__11), .D9_19(_RegFile_9__12), .D9_18(_RegFile_9__13),
		.D9_17(_RegFile_9__14), .D9_16(_RegFile_9__15), .D9_15(_RegFile_9__16),
		.D9_14(_RegFile_9__17), .D9_13(_RegFile_9__18), .D9_12(_RegFile_9__19),
		.D9_11(_RegFile_9__20), .D9_10(_RegFile_9__21), .D9_9(_RegFile_9__22),
		.D9_8(_RegFile_9__23), .D9_7(_RegFile_9__24), .D9_6(_RegFile_9__25),
		.D9_5(_RegFile_9__26), .D9_4(_RegFile_9__27), .D9_3(_RegFile_9__28),
		.D9_2(_RegFile_9__29), .D9_1(_RegFile_9__30), .D9_0(_RegFile_9__31),
		.D10_31(_RegFile_10__0), .D10_30(_RegFile_10__1), .D10_29(_RegFile_10__2),
		.D10_28(_RegFile_10__3), .D10_27(_RegFile_10__4), .D10_26(_RegFile_10__5),
		.D10_25(_RegFile_10__6), .D10_24(_RegFile_10__7), .D10_23(_RegFile_10__8),
		.D10_22(_RegFile_10__9), .D10_21(_RegFile_10__10), .D10_20(_RegFile_10__11),
		.D10_19(_RegFile_10__12), .D10_18(_RegFile_10__13), .D10_17(_RegFile_10__14),
		.D10_16(_RegFile_10__15), .D10_15(_RegFile_10__16), .D10_14(_RegFile_10__17),
		.D10_13(_RegFile_10__18), .D10_12(_RegFile_10__19), .D10_11(_RegFile_10__20),
		.D10_10(_RegFile_10__21), .D10_9(_RegFile_10__22), .D10_8(_RegFile_10__23),
		.D10_7(_RegFile_10__24), .D10_6(_RegFile_10__25), .D10_5(_RegFile_10__26),
		.D10_4(_RegFile_10__27), .D10_3(_RegFile_10__28), .D10_2(_RegFile_10__29),
		.D10_1(_RegFile_10__30), .D10_0(_RegFile_10__31), .D11_31(_RegFile_11__0),
		.D11_30(_RegFile_11__1), .D11_29(_RegFile_11__2), .D11_28(_RegFile_11__3),
		.D11_27(_RegFile_11__4), .D11_26(_RegFile_11__5), .D11_25(_RegFile_11__6),
		.D11_24(_RegFile_11__7), .D11_23(_RegFile_11__8), .D11_22(_RegFile_11__9),
		.D11_21(_RegFile_11__10), .D11_20(_RegFile_11__11), .D11_19(_RegFile_11__12),
		.D11_18(_RegFile_11__13), .D11_17(_RegFile_11__14), .D11_16(_RegFile_11__15),
		.D11_15(_RegFile_11__16), .D11_14(_RegFile_11__17), .D11_13(_RegFile_11__18),
		.D11_12(_RegFile_11__19), .D11_11(_RegFile_11__20), .D11_10(_RegFile_11__21),
		.D11_9(_RegFile_11__22), .D11_8(_RegFile_11__23), .D11_7(_RegFile_11__24),
		.D11_6(_RegFile_11__25), .D11_5(_RegFile_11__26), .D11_4(_RegFile_11__27),
		.D11_3(_RegFile_11__28), .D11_2(_RegFile_11__29), .D11_1(_RegFile_11__30),
		.D11_0(_RegFile_11__31), .D12_31(_RegFile_12__0), .D12_30(_RegFile_12__1),
		.D12_29(_RegFile_12__2), .D12_28(_RegFile_12__3), .D12_27(_RegFile_12__4),
		.D12_26(_RegFile_12__5), .D12_25(_RegFile_12__6), .D12_24(_RegFile_12__7),
		.D12_23(_RegFile_12__8), .D12_22(_RegFile_12__9), .D12_21(_RegFile_12__10),
		.D12_20(_RegFile_12__11), .D12_19(_RegFile_12__12), .D12_18(_RegFile_12__13),
		.D12_17(_RegFile_12__14), .D12_16(_RegFile_12__15), .D12_15(_RegFile_12__16),
		.D12_14(_RegFile_12__17), .D12_13(_RegFile_12__18), .D12_12(_RegFile_12__19),
		.D12_11(_RegFile_12__20), .D12_10(_RegFile_12__21), .D12_9(_RegFile_12__22),
		.D12_8(_RegFile_12__23), .D12_7(_RegFile_12__24), .D12_6(_RegFile_12__25),
		.D12_5(_RegFile_12__26), .D12_4(_RegFile_12__27), .D12_3(_RegFile_12__28),
		.D12_2(_RegFile_12__29), .D12_1(_RegFile_12__30), .D12_0(_RegFile_12__31),
		.D13_31(_RegFile_13__0), .D13_30(_RegFile_13__1), .D13_29(_RegFile_13__2),
		.D13_28(_RegFile_13__3), .D13_27(_RegFile_13__4), .D13_26(_RegFile_13__5),
		.D13_25(_RegFile_13__6), .D13_24(_RegFile_13__7), .D13_23(_RegFile_13__8),
		.D13_22(_RegFile_13__9), .D13_21(_RegFile_13__10), .D13_20(_RegFile_13__11),
		.D13_19(_RegFile_13__12), .D13_18(_RegFile_13__13), .D13_17(_RegFile_13__14),
		.D13_16(_RegFile_13__15), .D13_15(_RegFile_13__16), .D13_14(_RegFile_13__17),
		.D13_13(_RegFile_13__18), .D13_12(_RegFile_13__19), .D13_11(_RegFile_13__20),
		.D13_10(_RegFile_13__21), .D13_9(_RegFile_13__22), .D13_8(_RegFile_13__23),
		.D13_7(_RegFile_13__24), .D13_6(_RegFile_13__25), .D13_5(_RegFile_13__26),
		.D13_4(_RegFile_13__27), .D13_3(_RegFile_13__28), .D13_2(_RegFile_13__29),
		.D13_1(_RegFile_13__30), .D13_0(_RegFile_13__31), .D14_31(_RegFile_14__0),
		.D14_30(_RegFile_14__1), .D14_29(_RegFile_14__2), .D14_28(_RegFile_14__3),
		.D14_27(_RegFile_14__4), .D14_26(_RegFile_14__5), .D14_25(_RegFile_14__6),
		.D14_24(_RegFile_14__7), .D14_23(_RegFile_14__8), .D14_22(_RegFile_14__9),
		.D14_21(_RegFile_14__10), .D14_20(_RegFile_14__11), .D14_19(_RegFile_14__12),
		.D14_18(_RegFile_14__13), .D14_17(_RegFile_14__14), .D14_16(_RegFile_14__15),
		.D14_15(_RegFile_14__16), .D14_14(_RegFile_14__17), .D14_13(_RegFile_14__18),
		.D14_12(_RegFile_14__19), .D14_11(_RegFile_14__20), .D14_10(_RegFile_14__21),
		.D14_9(_RegFile_14__22), .D14_8(_RegFile_14__23), .D14_7(_RegFile_14__24),
		.D14_6(_RegFile_14__25), .D14_5(_RegFile_14__26), .D14_4(_RegFile_14__27),
		.D14_3(_RegFile_14__28), .D14_2(_RegFile_14__29), .D14_1(_RegFile_14__30),
		.D14_0(_RegFile_14__31), .D15_31(_RegFile_15__0), .D15_30(_RegFile_15__1),
		.D15_29(_RegFile_15__2), .D15_28(_RegFile_15__3), .D15_27(_RegFile_15__4),
		.D15_26(_RegFile_15__5), .D15_25(_RegFile_15__6), .D15_24(_RegFile_15__7),
		.D15_23(_RegFile_15__8), .D15_22(_RegFile_15__9), .D15_21(_RegFile_15__10),
		.D15_20(_RegFile_15__11), .D15_19(_RegFile_15__12), .D15_18(_RegFile_15__13),
		.D15_17(_RegFile_15__14), .D15_16(_RegFile_15__15), .D15_15(_RegFile_15__16),
		.D15_14(_RegFile_15__17), .D15_13(_RegFile_15__18), .D15_12(_RegFile_15__19),
		.D15_11(_RegFile_15__20), .D15_10(_RegFile_15__21), .D15_9(_RegFile_15__22),
		.D15_8(_RegFile_15__23), .D15_7(_RegFile_15__24), .D15_6(_RegFile_15__25),
		.D15_5(_RegFile_15__26), .D15_4(_RegFile_15__27), .D15_3(_RegFile_15__28),
		.D15_2(_RegFile_15__29), .D15_1(_RegFile_15__30), .D15_0(_RegFile_15__31),
		.D16_31(_RegFile_16__0), .D16_30(_RegFile_16__1), .D16_29(_RegFile_16__2),
		.D16_28(_RegFile_16__3), .D16_27(_RegFile_16__4), .D16_26(_RegFile_16__5),
		.D16_25(_RegFile_16__6), .D16_24(_RegFile_16__7), .D16_23(_RegFile_16__8),
		.D16_22(_RegFile_16__9), .D16_21(_RegFile_16__10), .D16_20(_RegFile_16__11),
		.D16_19(_RegFile_16__12), .D16_18(_RegFile_16__13), .D16_17(_RegFile_16__14),
		.D16_16(_RegFile_16__15), .D16_15(_RegFile_16__16), .D16_14(_RegFile_16__17),
		.D16_13(_RegFile_16__18), .D16_12(_RegFile_16__19), .D16_11(_RegFile_16__20),
		.D16_10(_RegFile_16__21), .D16_9(_RegFile_16__22), .D16_8(_RegFile_16__23),
		.D16_7(_RegFile_16__24), .D16_6(_RegFile_16__25), .D16_5(_RegFile_16__26),
		.D16_4(_RegFile_16__27), .D16_3(_RegFile_16__28), .D16_2(_RegFile_16__29),
		.D16_1(_RegFile_16__30), .D16_0(_RegFile_16__31), .D17_31(_RegFile_17__0),
		.D17_30(_RegFile_17__1), .D17_29(_RegFile_17__2), .D17_28(_RegFile_17__3),
		.D17_27(_RegFile_17__4), .D17_26(_RegFile_17__5), .D17_25(_RegFile_17__6),
		.D17_24(_RegFile_17__7), .D17_23(_RegFile_17__8), .D17_22(_RegFile_17__9),
		.D17_21(_RegFile_17__10), .D17_20(_RegFile_17__11), .D17_19(_RegFile_17__12),
		.D17_18(_RegFile_17__13), .D17_17(_RegFile_17__14), .D17_16(_RegFile_17__15),
		.D17_15(_RegFile_17__16), .D17_14(_RegFile_17__17), .D17_13(_RegFile_17__18),
		.D17_12(_RegFile_17__19), .D17_11(_RegFile_17__20), .D17_10(_RegFile_17__21),
		.D17_9(_RegFile_17__22), .D17_8(_RegFile_17__23), .D17_7(_RegFile_17__24),
		.D17_6(_RegFile_17__25), .D17_5(_RegFile_17__26), .D17_4(_RegFile_17__27),
		.D17_3(_RegFile_17__28), .D17_2(_RegFile_17__29), .D17_1(_RegFile_17__30),
		.D17_0(_RegFile_17__31), .D18_31(_RegFile_18__0), .D18_30(_RegFile_18__1),
		.D18_29(_RegFile_18__2), .D18_28(_RegFile_18__3), .D18_27(_RegFile_18__4),
		.D18_26(_RegFile_18__5), .D18_25(_RegFile_18__6), .D18_24(_RegFile_18__7),
		.D18_23(_RegFile_18__8), .D18_22(_RegFile_18__9), .D18_21(_RegFile_18__10),
		.D18_20(_RegFile_18__11), .D18_19(_RegFile_18__12), .D18_18(_RegFile_18__13),
		.D18_17(_RegFile_18__14), .D18_16(_RegFile_18__15), .D18_15(_RegFile_18__16),
		.D18_14(_RegFile_18__17), .D18_13(_RegFile_18__18), .D18_12(_RegFile_18__19),
		.D18_11(_RegFile_18__20), .D18_10(_RegFile_18__21), .D18_9(_RegFile_18__22),
		.D18_8(_RegFile_18__23), .D18_7(_RegFile_18__24), .D18_6(_RegFile_18__25),
		.D18_5(_RegFile_18__26), .D18_4(_RegFile_18__27), .D18_3(_RegFile_18__28),
		.D18_2(_RegFile_18__29), .D18_1(_RegFile_18__30), .D18_0(_RegFile_18__31),
		.D19_31(_RegFile_19__0), .D19_30(_RegFile_19__1), .D19_29(_RegFile_19__2),
		.D19_28(_RegFile_19__3), .D19_27(_RegFile_19__4), .D19_26(_RegFile_19__5),
		.D19_25(_RegFile_19__6), .D19_24(_RegFile_19__7), .D19_23(_RegFile_19__8),
		.D19_22(_RegFile_19__9), .D19_21(_RegFile_19__10), .D19_20(_RegFile_19__11),
		.D19_19(_RegFile_19__12), .D19_18(_RegFile_19__13), .D19_17(_RegFile_19__14),
		.D19_16(_RegFile_19__15), .D19_15(_RegFile_19__16), .D19_14(_RegFile_19__17),
		.D19_13(_RegFile_19__18), .D19_12(_RegFile_19__19), .D19_11(_RegFile_19__20),
		.D19_10(_RegFile_19__21), .D19_9(_RegFile_19__22), .D19_8(_RegFile_19__23),
		.D19_7(_RegFile_19__24), .D19_6(_RegFile_19__25), .D19_5(_RegFile_19__26),
		.D19_4(_RegFile_19__27), .D19_3(_RegFile_19__28), .D19_2(_RegFile_19__29),
		.D19_1(_RegFile_19__30), .D19_0(_RegFile_19__31), .D20_31(_RegFile_20__0),
		.D20_30(_RegFile_20__1), .D20_29(_RegFile_20__2), .D20_28(_RegFile_20__3),
		.D20_27(_RegFile_20__4), .D20_26(_RegFile_20__5), .D20_25(_RegFile_20__6),
		.D20_24(_RegFile_20__7), .D20_23(_RegFile_20__8), .D20_22(_RegFile_20__9),
		.D20_21(_RegFile_20__10), .D20_20(_RegFile_20__11), .D20_19(_RegFile_20__12),
		.D20_18(_RegFile_20__13), .D20_17(_RegFile_20__14), .D20_16(_RegFile_20__15),
		.D20_15(_RegFile_20__16), .D20_14(_RegFile_20__17), .D20_13(_RegFile_20__18),
		.D20_12(_RegFile_20__19), .D20_11(_RegFile_20__20), .D20_10(_RegFile_20__21),
		.D20_9(_RegFile_20__22), .D20_8(_RegFile_20__23), .D20_7(_RegFile_20__24),
		.D20_6(_RegFile_20__25), .D20_5(_RegFile_20__26), .D20_4(_RegFile_20__27),
		.D20_3(_RegFile_20__28), .D20_2(_RegFile_20__29), .D20_1(_RegFile_20__30),
		.D20_0(_RegFile_20__31), .D21_31(_RegFile_21__0), .D21_30(_RegFile_21__1),
		.D21_29(_RegFile_21__2), .D21_28(_RegFile_21__3), .D21_27(_RegFile_21__4),
		.D21_26(_RegFile_21__5), .D21_25(_RegFile_21__6), .D21_24(_RegFile_21__7),
		.D21_23(_RegFile_21__8), .D21_22(_RegFile_21__9), .D21_21(_RegFile_21__10),
		.D21_20(_RegFile_21__11), .D21_19(_RegFile_21__12), .D21_18(_RegFile_21__13),
		.D21_17(_RegFile_21__14), .D21_16(_RegFile_21__15), .D21_15(_RegFile_21__16),
		.D21_14(_RegFile_21__17), .D21_13(_RegFile_21__18), .D21_12(_RegFile_21__19),
		.D21_11(_RegFile_21__20), .D21_10(_RegFile_21__21), .D21_9(_RegFile_21__22),
		.D21_8(_RegFile_21__23), .D21_7(_RegFile_21__24), .D21_6(_RegFile_21__25),
		.D21_5(_RegFile_21__26), .D21_4(_RegFile_21__27), .D21_3(_RegFile_21__28),
		.D21_2(_RegFile_21__29), .D21_1(_RegFile_21__30), .D21_0(_RegFile_21__31),
		.D22_31(_RegFile_22__0), .D22_30(_RegFile_22__1), .D22_29(_RegFile_22__2),
		.D22_28(_RegFile_22__3), .D22_27(_RegFile_22__4), .D22_26(_RegFile_22__5),
		.D22_25(_RegFile_22__6), .D22_24(_RegFile_22__7), .D22_23(_RegFile_22__8),
		.D22_22(_RegFile_22__9), .D22_21(_RegFile_22__10), .D22_20(_RegFile_22__11),
		.D22_19(_RegFile_22__12), .D22_18(_RegFile_22__13), .D22_17(_RegFile_22__14),
		.D22_16(_RegFile_22__15), .D22_15(_RegFile_22__16), .D22_14(_RegFile_22__17),
		.D22_13(_RegFile_22__18), .D22_12(_RegFile_22__19), .D22_11(_RegFile_22__20),
		.D22_10(_RegFile_22__21), .D22_9(_RegFile_22__22), .D22_8(_RegFile_22__23),
		.D22_7(_RegFile_22__24), .D22_6(_RegFile_22__25), .D22_5(_RegFile_22__26),
		.D22_4(_RegFile_22__27), .D22_3(_RegFile_22__28), .D22_2(_RegFile_22__29),
		.D22_1(_RegFile_22__30), .D22_0(_RegFile_22__31), .D23_31(_RegFile_23__0),
		.D23_30(_RegFile_23__1), .D23_29(_RegFile_23__2), .D23_28(_RegFile_23__3),
		.D23_27(_RegFile_23__4), .D23_26(_RegFile_23__5), .D23_25(_RegFile_23__6),
		.D23_24(_RegFile_23__7), .D23_23(_RegFile_23__8), .D23_22(_RegFile_23__9),
		.D23_21(_RegFile_23__10), .D23_20(_RegFile_23__11), .D23_19(_RegFile_23__12),
		.D23_18(_RegFile_23__13), .D23_17(_RegFile_23__14), .D23_16(_RegFile_23__15),
		.D23_15(_RegFile_23__16), .D23_14(_RegFile_23__17), .D23_13(_RegFile_23__18),
		.D23_12(_RegFile_23__19), .D23_11(_RegFile_23__20), .D23_10(_RegFile_23__21),
		.D23_9(_RegFile_23__22), .D23_8(_RegFile_23__23), .D23_7(_RegFile_23__24),
		.D23_6(_RegFile_23__25), .D23_5(_RegFile_23__26), .D23_4(_RegFile_23__27),
		.D23_3(_RegFile_23__28), .D23_2(_RegFile_23__29), .D23_1(_RegFile_23__30),
		.D23_0(_RegFile_23__31), .D24_31(_RegFile_24__0), .D24_30(_RegFile_24__1),
		.D24_29(_RegFile_24__2), .D24_28(_RegFile_24__3), .D24_27(_RegFile_24__4),
		.D24_26(_RegFile_24__5), .D24_25(_RegFile_24__6), .D24_24(_RegFile_24__7),
		.D24_23(_RegFile_24__8), .D24_22(_RegFile_24__9), .D24_21(_RegFile_24__10),
		.D24_20(_RegFile_24__11), .D24_19(_RegFile_24__12), .D24_18(_RegFile_24__13),
		.D24_17(_RegFile_24__14), .D24_16(_RegFile_24__15), .D24_15(_RegFile_24__16),
		.D24_14(_RegFile_24__17), .D24_13(_RegFile_24__18), .D24_12(_RegFile_24__19),
		.D24_11(_RegFile_24__20), .D24_10(_RegFile_24__21), .D24_9(_RegFile_24__22),
		.D24_8(_RegFile_24__23), .D24_7(_RegFile_24__24), .D24_6(_RegFile_24__25),
		.D24_5(_RegFile_24__26), .D24_4(_RegFile_24__27), .D24_3(_RegFile_24__28),
		.D24_2(_RegFile_24__29), .D24_1(_RegFile_24__30), .D24_0(_RegFile_24__31),
		.D25_31(_RegFile_25__0), .D25_30(_RegFile_25__1), .D25_29(_RegFile_25__2),
		.D25_28(_RegFile_25__3), .D25_27(_RegFile_25__4), .D25_26(_RegFile_25__5),
		.D25_25(_RegFile_25__6), .D25_24(_RegFile_25__7), .D25_23(_RegFile_25__8),
		.D25_22(_RegFile_25__9), .D25_21(_RegFile_25__10), .D25_20(_RegFile_25__11),
		.D25_19(_RegFile_25__12), .D25_18(_RegFile_25__13), .D25_17(_RegFile_25__14),
		.D25_16(_RegFile_25__15), .D25_15(_RegFile_25__16), .D25_14(_RegFile_25__17),
		.D25_13(_RegFile_25__18), .D25_12(_RegFile_25__19), .D25_11(_RegFile_25__20),
		.D25_10(_RegFile_25__21), .D25_9(_RegFile_25__22), .D25_8(_RegFile_25__23),
		.D25_7(_RegFile_25__24), .D25_6(_RegFile_25__25), .D25_5(_RegFile_25__26),
		.D25_4(_RegFile_25__27), .D25_3(_RegFile_25__28), .D25_2(_RegFile_25__29),
		.D25_1(_RegFile_25__30), .D25_0(_RegFile_25__31), .D26_31(_RegFile_26__0),
		.D26_30(_RegFile_26__1), .D26_29(_RegFile_26__2), .D26_28(_RegFile_26__3),
		.D26_27(_RegFile_26__4), .D26_26(_RegFile_26__5), .D26_25(_RegFile_26__6),
		.D26_24(_RegFile_26__7), .D26_23(_RegFile_26__8), .D26_22(_RegFile_26__9),
		.D26_21(_RegFile_26__10), .D26_20(_RegFile_26__11), .D26_19(_RegFile_26__12),
		.D26_18(_RegFile_26__13), .D26_17(_RegFile_26__14), .D26_16(_RegFile_26__15),
		.D26_15(_RegFile_26__16), .D26_14(_RegFile_26__17), .D26_13(_RegFile_26__18),
		.D26_12(_RegFile_26__19), .D26_11(_RegFile_26__20), .D26_10(_RegFile_26__21),
		.D26_9(_RegFile_26__22), .D26_8(_RegFile_26__23), .D26_7(_RegFile_26__24),
		.D26_6(_RegFile_26__25), .D26_5(_RegFile_26__26), .D26_4(_RegFile_26__27),
		.D26_3(_RegFile_26__28), .D26_2(_RegFile_26__29), .D26_1(_RegFile_26__30),
		.D26_0(_RegFile_26__31), .D27_31(_RegFile_27__0), .D27_30(_RegFile_27__1),
		.D27_29(_RegFile_27__2), .D27_28(_RegFile_27__3), .D27_27(_RegFile_27__4),
		.D27_26(_RegFile_27__5), .D27_25(_RegFile_27__6), .D27_24(_RegFile_27__7),
		.D27_23(_RegFile_27__8), .D27_22(_RegFile_27__9), .D27_21(_RegFile_27__10),
		.D27_20(_RegFile_27__11), .D27_19(_RegFile_27__12), .D27_18(_RegFile_27__13),
		.D27_17(_RegFile_27__14), .D27_16(_RegFile_27__15), .D27_15(_RegFile_27__16),
		.D27_14(_RegFile_27__17), .D27_13(_RegFile_27__18), .D27_12(_RegFile_27__19),
		.D27_11(_RegFile_27__20), .D27_10(_RegFile_27__21), .D27_9(_RegFile_27__22),
		.D27_8(_RegFile_27__23), .D27_7(_RegFile_27__24), .D27_6(_RegFile_27__25),
		.D27_5(_RegFile_27__26), .D27_4(_RegFile_27__27), .D27_3(_RegFile_27__28),
		.D27_2(_RegFile_27__29), .D27_1(_RegFile_27__30), .D27_0(_RegFile_27__31),
		.D28_31(_RegFile_28__0), .D28_30(_RegFile_28__1), .D28_29(_RegFile_28__2),
		.D28_28(_RegFile_28__3), .D28_27(_RegFile_28__4), .D28_26(_RegFile_28__5),
		.D28_25(_RegFile_28__6), .D28_24(_RegFile_28__7), .D28_23(_RegFile_28__8),
		.D28_22(_RegFile_28__9), .D28_21(_RegFile_28__10), .D28_20(_RegFile_28__11),
		.D28_19(_RegFile_28__12), .D28_18(_RegFile_28__13), .D28_17(_RegFile_28__14),
		.D28_16(_RegFile_28__15), .D28_15(_RegFile_28__16), .D28_14(_RegFile_28__17),
		.D28_13(_RegFile_28__18), .D28_12(_RegFile_28__19), .D28_11(_RegFile_28__20),
		.D28_10(_RegFile_28__21), .D28_9(_RegFile_28__22), .D28_8(_RegFile_28__23),
		.D28_7(_RegFile_28__24), .D28_6(_RegFile_28__25), .D28_5(_RegFile_28__26),
		.D28_4(_RegFile_28__27), .D28_3(_RegFile_28__28), .D28_2(_RegFile_28__29),
		.D28_1(_RegFile_28__30), .D28_0(_RegFile_28__31), .D29_31(_RegFile_29__0),
		.D29_30(_RegFile_29__1), .D29_29(_RegFile_29__2), .D29_28(_RegFile_29__3),
		.D29_27(_RegFile_29__4), .D29_26(_RegFile_29__5), .D29_25(_RegFile_29__6),
		.D29_24(_RegFile_29__7), .D29_23(_RegFile_29__8), .D29_22(_RegFile_29__9),
		.D29_21(_RegFile_29__10), .D29_20(_RegFile_29__11), .D29_19(_RegFile_29__12),
		.D29_18(_RegFile_29__13), .D29_17(_RegFile_29__14), .D29_16(_RegFile_29__15),
		.D29_15(_RegFile_29__16), .D29_14(_RegFile_29__17), .D29_13(_RegFile_29__18),
		.D29_12(_RegFile_29__19), .D29_11(_RegFile_29__20), .D29_10(_RegFile_29__21),
		.D29_9(_RegFile_29__22), .D29_8(_RegFile_29__23), .D29_7(_RegFile_29__24),
		.D29_6(_RegFile_29__25), .D29_5(_RegFile_29__26), .D29_4(_RegFile_29__27),
		.D29_3(_RegFile_29__28), .D29_2(_RegFile_29__29), .D29_1(_RegFile_29__30),
		.D29_0(_RegFile_29__31), .D30_31(_RegFile_30__0), .D30_30(_RegFile_30__1),
		.D30_29(_RegFile_30__2), .D30_28(_RegFile_30__3), .D30_27(_RegFile_30__4),
		.D30_26(_RegFile_30__5), .D30_25(_RegFile_30__6), .D30_24(_RegFile_30__7),
		.D30_23(_RegFile_30__8), .D30_22(_RegFile_30__9), .D30_21(_RegFile_30__10),
		.D30_20(_RegFile_30__11), .D30_19(_RegFile_30__12), .D30_18(_RegFile_30__13),
		.D30_17(_RegFile_30__14), .D30_16(_RegFile_30__15), .D30_15(_RegFile_30__16),
		.D30_14(_RegFile_30__17), .D30_13(_RegFile_30__18), .D30_12(_RegFile_30__19),
		.D30_11(_RegFile_30__20), .D30_10(_RegFile_30__21), .D30_9(_RegFile_30__22),
		.D30_8(_RegFile_30__23), .D30_7(_RegFile_30__24), .D30_6(_RegFile_30__25),
		.D30_5(_RegFile_30__26), .D30_4(_RegFile_30__27), .D30_3(_RegFile_30__28),
		.D30_2(_RegFile_30__29), .D30_1(_RegFile_30__30), .D30_0(_RegFile_30__31),
		.D31_31(_RegFile_31__0), .D31_30(_RegFile_31__1), .D31_29(_RegFile_31__2),
		.D31_28(_RegFile_31__3), .D31_27(_RegFile_31__4), .D31_26(_RegFile_31__5),
		.D31_25(_RegFile_31__6), .D31_24(_RegFile_31__7), .D31_23(_RegFile_31__8),
		.D31_22(_RegFile_31__9), .D31_21(_RegFile_31__10), .D31_20(_RegFile_31__11),
		.D31_19(_RegFile_31__12), .D31_18(_RegFile_31__13), .D31_17(_RegFile_31__14),
		.D31_16(_RegFile_31__15), .D31_15(_RegFile_31__16), .D31_14(_RegFile_31__17),
		.D31_13(_RegFile_31__18), .D31_12(_RegFile_31__19), .D31_11(_RegFile_31__20),
		.D31_10(_RegFile_31__21), .D31_9(_RegFile_31__22), .D31_8(_RegFile_31__23),
		.D31_7(_RegFile_31__24), .D31_6(_RegFile_31__25), .D31_5(_RegFile_31__26),
		.D31_4(_RegFile_31__27), .D31_3(_RegFile_31__28), .D31_2(_RegFile_31__29),
		.D31_1(_RegFile_31__30), .D31_0(_RegFile_31__31), .S0(n857), .S1(n339),
		.S2(n848), .S3(n337), .S4(n802), .Z_31(N535), .Z_30(N534), .Z_29(N533),
		.Z_28(N532), .Z_27(N531), .Z_26(N530), .Z_25(N529), .Z_24(N528), .Z_23(N527),
		.Z_22(N526), .Z_21(N525), .Z_20(N524), .Z_19(N523), .Z_18(N522), .Z_17(N521),
		.Z_16(N520), .Z_15(N519), .Z_14(N518), .Z_13(N517), .Z_12(N516), .Z_11(N515),
		.Z_10(N514), .Z_9(N513), .Z_8(N512), .Z_7(N511), .Z_6(N510), .Z_5(N509),
		.Z_4(N508), .Z_3(N507), .Z_2(N506), .Z_1(N505), .Z_0(N504) );
	smlatnr_1 CLI_reg__master ( .q(CLI_reg__m2s), .qb(), .d(n2641), .sdi(test_si),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 CLI_reg__slave ( .q(CLI), .qb(n4386), .d(CLI_reg__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_0__master ( .q(Cause_Reg_reg_0__m2s), .qb(), .d(n2642),
		.sdi(n4386), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_0__slave ( .q(Cause_Reg_0), .qb(n627), .d(Cause_Reg_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_10__master ( .q(Cause_Reg_reg_10__m2s), .qb(),
		.d(n2652), .sdi(n618), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_10__slave ( .q(Cause_Reg_10), .qb(n617), .d(Cause_Reg_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_11__master ( .q(Cause_Reg_reg_11__m2s), .qb(),
		.d(n2653), .sdi(n617), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_11__slave ( .q(Cause_Reg_11), .qb(n616), .d(Cause_Reg_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_12__master ( .q(Cause_Reg_reg_12__m2s), .qb(),
		.d(n2654), .sdi(n616), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_12__slave ( .q(Cause_Reg_12), .qb(n615), .d(Cause_Reg_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_13__master ( .q(Cause_Reg_reg_13__m2s), .qb(),
		.d(n2655), .sdi(n615), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_13__slave ( .q(Cause_Reg_13), .qb(n614), .d(Cause_Reg_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_14__master ( .q(Cause_Reg_reg_14__m2s), .qb(),
		.d(n2656), .sdi(n614), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_14__slave ( .q(Cause_Reg_14), .qb(n613), .d(Cause_Reg_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_15__master ( .q(Cause_Reg_reg_15__m2s), .qb(),
		.d(n2657), .sdi(n613), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_15__slave ( .q(Cause_Reg_15), .qb(n612), .d(Cause_Reg_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_16__master ( .q(Cause_Reg_reg_16__m2s), .qb(),
		.d(n2658), .sdi(n612), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_16__slave ( .q(Cause_Reg_16), .qb(n611), .d(Cause_Reg_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_17__master ( .q(Cause_Reg_reg_17__m2s), .qb(),
		.d(n2659), .sdi(n611), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_17__slave ( .q(Cause_Reg_17), .qb(n610), .d(Cause_Reg_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_18__master ( .q(Cause_Reg_reg_18__m2s), .qb(),
		.d(n2660), .sdi(n610), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_18__slave ( .q(Cause_Reg_18), .qb(n609), .d(Cause_Reg_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_19__master ( .q(Cause_Reg_reg_19__m2s), .qb(),
		.d(n2661), .sdi(n609), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_19__slave ( .q(Cause_Reg_19), .qb(n608), .d(Cause_Reg_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_1__master ( .q(Cause_Reg_reg_1__m2s), .qb(), .d(n2643),
		.sdi(n627), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_1__slave ( .q(Cause_Reg_1), .qb(n626), .d(Cause_Reg_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_20__master ( .q(Cause_Reg_reg_20__m2s), .qb(),
		.d(n2662), .sdi(n608), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_20__slave ( .q(Cause_Reg_20), .qb(n607), .d(Cause_Reg_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_21__master ( .q(Cause_Reg_reg_21__m2s), .qb(),
		.d(n2663), .sdi(n607), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_21__slave ( .q(Cause_Reg_21), .qb(n606), .d(Cause_Reg_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_22__master ( .q(Cause_Reg_reg_22__m2s), .qb(),
		.d(n2664), .sdi(n606), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_22__slave ( .q(Cause_Reg_22), .qb(n605), .d(Cause_Reg_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_23__master ( .q(Cause_Reg_reg_23__m2s), .qb(),
		.d(n2665), .sdi(n605), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_23__slave ( .q(Cause_Reg_23), .qb(n604), .d(Cause_Reg_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_24__master ( .q(Cause_Reg_reg_24__m2s), .qb(),
		.d(n2666), .sdi(n604), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_24__slave ( .q(Cause_Reg_24), .qb(n603), .d(Cause_Reg_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_25__master ( .q(Cause_Reg_reg_25__m2s), .qb(),
		.d(n2667), .sdi(n603), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_25__slave ( .q(Cause_Reg_25), .qb(n602), .d(Cause_Reg_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_26__master ( .q(Cause_Reg_reg_26__m2s), .qb(),
		.d(n2668), .sdi(n602), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_26__slave ( .q(Cause_Reg_26), .qb(n601), .d(Cause_Reg_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_27__master ( .q(Cause_Reg_reg_27__m2s), .qb(),
		.d(n2669), .sdi(n601), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_27__slave ( .q(Cause_Reg_27), .qb(n600), .d(Cause_Reg_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_28__master ( .q(Cause_Reg_reg_28__m2s), .qb(),
		.d(n2670), .sdi(n600), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_28__slave ( .q(Cause_Reg_28), .qb(n599), .d(Cause_Reg_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_29__master ( .q(Cause_Reg_reg_29__m2s), .qb(),
		.d(n2671), .sdi(n599), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_29__slave ( .q(Cause_Reg_29), .qb(n598), .d(Cause_Reg_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_2__master ( .q(Cause_Reg_reg_2__m2s), .qb(), .d(n2644),
		.sdi(n626), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n953), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_2__slave ( .q(Cause_Reg_2), .qb(n625), .d(Cause_Reg_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n953), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_30__master ( .q(Cause_Reg_reg_30__m2s), .qb(),
		.d(n2672), .sdi(n598), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_30__slave ( .q(Cause_Reg_30), .qb(n597), .d(Cause_Reg_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_31__master ( .q(Cause_Reg_reg_31__m2s), .qb(),
		.d(n2673), .sdi(n597), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_31__slave ( .q(Cause_Reg_31), .qb(n596), .d(Cause_Reg_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_3__master ( .q(Cause_Reg_reg_3__m2s), .qb(), .d(n2645),
		.sdi(n625), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_3__slave ( .q(Cause_Reg_3), .qb(n624), .d(Cause_Reg_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_4__master ( .q(Cause_Reg_reg_4__m2s), .qb(), .d(n2646),
		.sdi(n624), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_4__slave ( .q(Cause_Reg_4), .qb(n623), .d(Cause_Reg_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_5__master ( .q(Cause_Reg_reg_5__m2s), .qb(), .d(n2647),
		.sdi(n623), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_5__slave ( .q(Cause_Reg_5), .qb(n622), .d(Cause_Reg_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_6__master ( .q(Cause_Reg_reg_6__m2s), .qb(), .d(n2648),
		.sdi(n622), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_6__slave ( .q(Cause_Reg_6), .qb(n621), .d(Cause_Reg_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_7__master ( .q(Cause_Reg_reg_7__m2s), .qb(), .d(n2649),
		.sdi(n621), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_7__slave ( .q(Cause_Reg_7), .qb(n620), .d(Cause_Reg_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_8__master ( .q(Cause_Reg_reg_8__m2s), .qb(), .d(n2650),
		.sdi(n620), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_8__slave ( .q(Cause_Reg_8), .qb(n619), .d(Cause_Reg_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Cause_Reg_reg_9__master ( .q(Cause_Reg_reg_9__m2s), .qb(), .d(n2651),
		.sdi(n619), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 Cause_Reg_reg_9__slave ( .q(Cause_Reg_9), .qb(n618), .d(Cause_Reg_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_0__master ( .q(EPC_reg_0__m2s), .qb(), .d(n2674), .sdi(n596),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_0__slave ( .q(EPC_0), .qb(n595), .d(EPC_reg_0__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_10__master ( .q(EPC_reg_10__m2s), .qb(), .d(n2684), .sdi(EPC_9),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_10__slave ( .q(EPC_10), .qb(n593), .d(EPC_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_11__master ( .q(EPC_reg_11__m2s), .qb(), .d(n2685), .sdi(EPC_10),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_11__slave ( .q(EPC_11), .qb(n592), .d(EPC_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_12__master ( .q(EPC_reg_12__m2s), .qb(), .d(n2686), .sdi(EPC_11),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_12__slave ( .q(EPC_12), .qb(n591), .d(EPC_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_13__master ( .q(EPC_reg_13__m2s), .qb(), .d(n2687), .sdi(EPC_12),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_13__slave ( .q(EPC_13), .qb(n590), .d(EPC_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_14__master ( .q(EPC_reg_14__m2s), .qb(), .d(n2688), .sdi(EPC_13),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_14__slave ( .q(EPC_14), .qb(n589), .d(EPC_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_15__master ( .q(EPC_reg_15__m2s), .qb(), .d(n2689), .sdi(EPC_14),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_15__slave ( .q(EPC_15), .qb(n588), .d(EPC_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_16__master ( .q(EPC_reg_16__m2s), .qb(), .d(n2690), .sdi(n588),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_16__slave ( .q(EPC_16), .qb(n587), .d(EPC_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_17__master ( .q(EPC_reg_17__m2s), .qb(), .d(n2691), .sdi(EPC_16),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_17__slave ( .q(EPC_17), .qb(n586), .d(EPC_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_18__master ( .q(EPC_reg_18__m2s), .qb(), .d(n2692), .sdi(EPC_17),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_18__slave ( .q(EPC_18), .qb(n585), .d(EPC_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_19__master ( .q(EPC_reg_19__m2s), .qb(), .d(n2693), .sdi(EPC_18),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_19__slave ( .q(EPC_19), .qb(n584), .d(EPC_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_1__master ( .q(EPC_reg_1__m2s), .qb(), .d(n2675), .sdi(EPC_0),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n952), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_1__slave ( .q(EPC_1), .qb(n594), .d(EPC_reg_1__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n952), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_20__master ( .q(EPC_reg_20__m2s), .qb(), .d(n2694), .sdi(EPC_19),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_20__slave ( .q(EPC_20), .qb(n583), .d(EPC_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_21__master ( .q(EPC_reg_21__m2s), .qb(), .d(n2695), .sdi(EPC_20),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_21__slave ( .q(EPC_21), .qb(n4383), .d(EPC_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_22__master ( .q(EPC_reg_22__m2s), .qb(), .d(n2696), .sdi(n4383),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_22__slave ( .q(EPC_22), .qb(n4382), .d(EPC_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_23__master ( .q(EPC_reg_23__m2s), .qb(), .d(n2697), .sdi(n4382),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_23__slave ( .q(EPC_23), .qb(n4381), .d(EPC_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_24__master ( .q(EPC_reg_24__m2s), .qb(), .d(n2698), .sdi(n4381),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_24__slave ( .q(EPC_24), .qb(n4380), .d(EPC_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_25__master ( .q(EPC_reg_25__m2s), .qb(), .d(n2699), .sdi(n4380),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_25__slave ( .q(EPC_25), .qb(n4379), .d(EPC_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_26__master ( .q(EPC_reg_26__m2s), .qb(), .d(n2700), .sdi(n4379),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_26__slave ( .q(EPC_26), .qb(n582), .d(EPC_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_27__master ( .q(EPC_reg_27__m2s), .qb(), .d(n2701), .sdi(n582),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_27__slave ( .q(EPC_27), .qb(n581), .d(EPC_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_28__master ( .q(EPC_reg_28__m2s), .qb(), .d(n2702), .sdi(n581),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_28__slave ( .q(EPC_28), .qb(n580), .d(EPC_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_29__master ( .q(EPC_reg_29__m2s), .qb(), .d(n2703), .sdi(n580),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_29__slave ( .q(EPC_29), .qb(n579), .d(EPC_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_2__master ( .q(EPC_reg_2__m2s), .qb(), .d(n2676), .sdi(EPC_1),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n954), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_2__slave ( .q(EPC_2), .qb(n4385), .d(EPC_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n954), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_30__master ( .q(EPC_reg_30__m2s), .qb(), .d(n2704), .sdi(n579),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_30__slave ( .q(EPC_30), .qb(n662), .d(EPC_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_31__master ( .q(EPC_reg_31__m2s), .qb(), .d(_EPC_reg_31_net69891),
		.sdi(EPC_30), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_31__slave ( .q(EPC_31), .qb(n578), .d(EPC_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_3__master ( .q(EPC_reg_3__m2s), .qb(), .d(n2677), .sdi(n4385),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_3__slave ( .q(EPC_3), .qb(n4384), .d(EPC_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_4__master ( .q(EPC_reg_4__m2s), .qb(), .d(n2678), .sdi(n4384),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_4__slave ( .q(EPC_4), .qb(n577), .d(EPC_reg_4__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_5__master ( .q(EPC_reg_5__m2s), .qb(), .d(n2679), .sdi(EPC_4),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_5__slave ( .q(EPC_5), .qb(n576), .d(EPC_reg_5__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_6__master ( .q(EPC_reg_6__m2s), .qb(), .d(n2680), .sdi(EPC_5),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_6__slave ( .q(EPC_6), .qb(n575), .d(EPC_reg_6__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_7__master ( .q(EPC_reg_7__m2s), .qb(), .d(n2681), .sdi(EPC_6),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_7__slave ( .q(EPC_7), .qb(n574), .d(EPC_reg_7__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_8__master ( .q(EPC_reg_8__m2s), .qb(), .d(n2682), .sdi(EPC_7),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_8__slave ( .q(EPC_8), .qb(n573), .d(EPC_reg_8__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 EPC_reg_9__master ( .q(EPC_reg_9__m2s), .qb(), .d(n2683), .sdi(EPC_8),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 EPC_reg_9__slave ( .q(EPC_9), .qb(n572), .d(EPC_reg_9__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_function_field_reg_0__master ( .q(IR_function_field_reg_0__m2s),
		.qb(), .d(n3764), .sdi(EPC_31), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n955), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_function_field_reg_0__slave ( .q(IR_function_field[0]), .qb(n1859),
		.d(IR_function_field_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_function_field_reg_1__master ( .q(IR_function_field_reg_1__m2s),
		.qb(), .d(n3765), .sdi(n1859), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_function_field_reg_1__slave ( .q(IR_function_field[1]), .qb(n1860),
		.d(IR_function_field_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_function_field_reg_2__master ( .q(IR_function_field_reg_2__m2s),
		.qb(), .d(n3766), .sdi(n1860), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_function_field_reg_2__slave ( .q(IR_function_field[2]), .qb(n1861),
		.d(IR_function_field_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_function_field_reg_3__master ( .q(IR_function_field_reg_3__m2s),
		.qb(), .d(n3767), .sdi(n1861), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_function_field_reg_3__slave ( .q(IR_function_field[3]), .qb(n1862),
		.d(IR_function_field_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_function_field_reg_4__master ( .q(IR_function_field_reg_4__m2s),
		.qb(), .d(n3768), .sdi(n1862), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_function_field_reg_4__slave ( .q(IR_function_field[4]), .qb(n1863),
		.d(IR_function_field_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_function_field_reg_5__master ( .q(IR_function_field_reg_5__m2s),
		.qb(), .d(n3769), .sdi(n1863), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_function_field_reg_5__slave ( .q(IR_function_field[5]), .qb(n4378),
		.d(IR_function_field_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_opcode_field_reg_0__master ( .q(IR_opcode_field_reg_0__m2s),
		.qb(), .d(n3770), .sdi(n4378), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 IR_opcode_field_reg_0__slave ( .q(n4454), .qb(n4377), .d(IR_opcode_field_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_opcode_field_reg_1__master ( .q(IR_opcode_field_reg_1__m2s),
		.qb(), .d(n3771), .sdi(n4377), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 IR_opcode_field_reg_1__slave ( .q(n4453), .qb(n4376), .d(IR_opcode_field_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_opcode_field_reg_2__master ( .q(IR_opcode_field_reg_2__m2s),
		.qb(), .d(n3772), .sdi(n4376), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 IR_opcode_field_reg_2__slave ( .q(n4452), .qb(n4375), .d(IR_opcode_field_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_opcode_field_reg_3__master ( .q(IR_opcode_field_reg_3__m2s),
		.qb(), .d(n3773), .sdi(n4375), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 IR_opcode_field_reg_3__slave ( .q(IR_opcode_field[3]), .qb(n4374),
		.d(IR_opcode_field_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_opcode_field_reg_4__master ( .q(IR_opcode_field_reg_4__m2s),
		.qb(), .d(n3774), .sdi(n4374), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 IR_opcode_field_reg_4__slave ( .q(IR_opcode_field[4]), .qb(n4373),
		.d(IR_opcode_field_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 IR_opcode_field_reg_5__master ( .q(IR_opcode_field_reg_5__m2s),
		.qb(), .d(n3775), .sdi(n4373), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 IR_opcode_field_reg_5__slave ( .q(IR_opcode_field[5]), .qb(n4372),
		.d(IR_opcode_field_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_0__master ( .q(Imm_reg_0__m2s), .qb(), .d(n3791), .sdi(n4372),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_0__slave ( .q(N6328), .qb(n813), .d(Imm_reg_0__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_10__master ( .q(Imm_reg_10__m2s), .qb(), .d(n3801), .sdi(n873),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_10__slave ( .q(N6348), .qb(n4371), .d(Imm_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_11__master ( .q(Imm_reg_11__m2s), .qb(), .d(n3802), .sdi(n4371),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_11__slave ( .q(N6350), .qb(n786), .d(Imm_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_12__master ( .q(Imm_reg_12__m2s), .qb(), .d(n3803), .sdi(n786),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_12__slave ( .q(N6352), .qb(n779), .d(Imm_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_13__master ( .q(Imm_reg_13__m2s), .qb(), .d(n3804), .sdi(n779),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_13__slave ( .q(N6354), .qb(n4370), .d(Imm_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_14__master ( .q(Imm_reg_14__m2s), .qb(), .d(n3805), .sdi(n4370),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_14__slave ( .q(N6356), .qb(n647), .d(Imm_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_15__master ( .q(Imm_reg_15__m2s), .qb(), .d(n3806), .sdi(n647),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_15__slave ( .q(N6358), .qb(n829), .d(Imm_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_16__master ( .q(Imm_reg_16__m2s), .qb(), .d(n3807), .sdi(n829),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_16__slave ( .q(N6360), .qb(n648), .d(Imm_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_17__master ( .q(Imm_reg_17__m2s), .qb(), .d(n3808), .sdi(n648),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_17__slave ( .q(N6362), .qb(n803), .d(Imm_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_18__master ( .q(Imm_reg_18__m2s), .qb(), .d(n3809), .sdi(n803),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_18__slave ( .q(N6364), .qb(n778), .d(Imm_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_19__master ( .q(Imm_reg_19__m2s), .qb(), .d(n3810), .sdi(n778),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_19__slave ( .q(N6366), .qb(n775), .d(Imm_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_1__master ( .q(Imm_reg_1__m2s), .qb(), .d(n3792), .sdi(n813),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_1__slave ( .q(Imm[1]), .qb(n720), .d(Imm_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_20__master ( .q(Imm_reg_20__m2s), .qb(), .d(n3811), .sdi(n775),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_20__slave ( .q(N6368), .qb(n732), .d(Imm_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_21__master ( .q(Imm_reg_21__m2s), .qb(), .d(n3812), .sdi(n732),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_21__slave ( .q(N6370), .qb(n649), .d(Imm_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_22__master ( .q(Imm_reg_22__m2s), .qb(), .d(n3813), .sdi(n649),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_22__slave ( .q(Imm[22]), .qb(n789), .d(Imm_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_23__master ( .q(Imm_reg_23__m2s), .qb(), .d(n3814), .sdi(n789),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_23__slave ( .q(Imm[23]), .qb(n827), .d(Imm_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_24__master ( .q(Imm_reg_24__m2s), .qb(), .d(n3815), .sdi(n827),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_24__slave ( .q(N6376), .qb(n654), .d(Imm_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_25__master ( .q(Imm_reg_25__m2s), .qb(), .d(n3816), .sdi(n654),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n951), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_25__slave ( .q(Imm[25]), .qb(n816), .d(Imm_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n951), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_26__master ( .q(Imm_reg_26__m2s), .qb(), .d(n3817), .sdi(n816),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_26__slave ( .q(N6380), .qb(n735), .d(Imm_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_27__master ( .q(Imm_reg_27__m2s), .qb(), .d(n3818), .sdi(n735),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_27__slave ( .q(N6382), .qb(n765), .d(Imm_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_28__master ( .q(Imm_reg_28__m2s), .qb(), .d(n3819), .sdi(n765),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_28__slave ( .q(N6384), .qb(n696), .d(Imm_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_29__master ( .q(Imm_reg_29__m2s), .qb(), .d(n3820), .sdi(n696),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_29__slave ( .q(N6386), .qb(n762), .d(Imm_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_2__master ( .q(Imm_reg_2__m2s), .qb(), .d(n3793), .sdi(n720),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_2__slave ( .q(N6332), .qb(n870), .d(Imm_reg_2__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_30__master ( .q(Imm_reg_30__m2s), .qb(), .d(n3821), .sdi(n762),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_30__slave ( .q(N6388), .qb(n701), .d(Imm_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_31__master ( .q(Imm_reg_31__m2s), .qb(), .d(n3822), .sdi(n701),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_31__slave ( .q(N6390), .qb(n4369), .d(Imm_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_3__master ( .q(Imm_reg_3__m2s), .qb(), .d(n3794), .sdi(n870),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_3__slave ( .q(N6334), .qb(n886), .d(Imm_reg_3__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_4__master ( .q(Imm_reg_4__m2s), .qb(), .d(n3795), .sdi(n886),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_4__slave ( .q(N6336), .qb(n871), .d(Imm_reg_4__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_5__master ( .q(Imm_reg_5__m2s), .qb(), .d(n3796), .sdi(n871),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_5__slave ( .q(N6338), .qb(n845), .d(Imm_reg_5__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_6__master ( .q(Imm_reg_6__m2s), .qb(), .d(n3797), .sdi(n845),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_6__slave ( .q(N6340), .qb(n643), .d(Imm_reg_6__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_7__master ( .q(Imm_reg_7__m2s), .qb(), .d(n3798), .sdi(n643),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_7__slave ( .q(N6342), .qb(n734), .d(Imm_reg_7__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_8__master ( .q(Imm_reg_8__m2s), .qb(), .d(n3799), .sdi(n734),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 Imm_reg_8__slave ( .q(N6344), .qb(n872), .d(Imm_reg_8__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 Imm_reg_9__master ( .q(Imm_reg_9__m2s), .qb(), .d(n3800), .sdi(n872),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 Imm_reg_9__slave ( .q(N6346), .qb(n873), .d(Imm_reg_9__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	inv_2 U10 ( .x(n554), .a(n1547) );
	inv_2 U100 ( .x(n1382), .a(N449) );
	or2_2 U1000 ( .x(n1767), .a(n3936), .b(n3940) );
	mux2_2 U1001 ( .x(n3285), .d0(_RegFile_13__0), .sl(n1830), .d1(WB_data[0]) );
	mux2_2 U1002 ( .x(n3286), .d0(_RegFile_13__1), .sl(n1830), .d1(WB_data[1]) );
	mux2_2 U1003 ( .x(n3287), .d0(_RegFile_13__2), .sl(n1830), .d1(WB_data[2]) );
	mux2_2 U1004 ( .x(n3288), .d0(_RegFile_13__3), .sl(n1830), .d1(WB_data[3]) );
	mux2_2 U1005 ( .x(n3289), .d0(_RegFile_13__4), .sl(n1830), .d1(WB_data[4]) );
	mux2_2 U1006 ( .x(n3290), .d0(_RegFile_13__5), .sl(n1830), .d1(WB_data[5]) );
	mux2_2 U1007 ( .x(n3291), .d0(_RegFile_13__6), .sl(n1830), .d1(WB_data[6]) );
	mux2_2 U1008 ( .x(n3292), .d0(_RegFile_13__7), .sl(n1830), .d1(WB_data[7]) );
	mux2i_1 U1009 ( .x(n3294), .d0(n1983), .sl(n1830), .d1(n1801) );
	inv_2 U101 ( .x(n1399), .a(N456) );
	mux2i_1 U1010 ( .x(n3295), .d0(n1960), .sl(n1830), .d1(n1778) );
	mux2i_1 U1011 ( .x(n3296), .d0(n1961), .sl(n1830), .d1(n1779) );
	mux2i_1 U1012 ( .x(n3297), .d0(n1962), .sl(n1830), .d1(n1780) );
	mux2i_1 U1013 ( .x(n3298), .d0(n1963), .sl(n1830), .d1(n1781) );
	mux2i_1 U1014 ( .x(n3299), .d0(n1964), .sl(n1830), .d1(n1782) );
	mux2i_1 U1015 ( .x(n3300), .d0(n1965), .sl(n1830), .d1(n1783) );
	mux2i_1 U1016 ( .x(n3301), .d0(n1966), .sl(n1830), .d1(n1784) );
	mux2i_1 U1017 ( .x(n3302), .d0(n1967), .sl(n1830), .d1(n1785) );
	mux2i_1 U1018 ( .x(n3303), .d0(n1968), .sl(n1830), .d1(n1786) );
	mux2i_1 U1019 ( .x(n3304), .d0(n1969), .sl(n1830), .d1(n1787) );
	nand2i_2 U102 ( .x(n1520), .a(n1515), .b(n1521) );
	mux2i_1 U1020 ( .x(n3305), .d0(n1970), .sl(n1830), .d1(n1788) );
	mux2i_1 U1021 ( .x(n3306), .d0(n1971), .sl(n1830), .d1(n1789) );
	mux2i_1 U1022 ( .x(n3307), .d0(n1972), .sl(n1830), .d1(n1790) );
	mux2i_1 U1023 ( .x(n3308), .d0(n1973), .sl(n1830), .d1(n1791) );
	mux2i_1 U1024 ( .x(n3309), .d0(n1974), .sl(n1830), .d1(n1792) );
	mux2i_1 U1025 ( .x(n3310), .d0(n1975), .sl(n1830), .d1(n1793) );
	mux2i_1 U1026 ( .x(n3311), .d0(n1976), .sl(n1830), .d1(n1794) );
	mux2i_1 U1027 ( .x(n3312), .d0(n1977), .sl(n1830), .d1(n1795) );
	mux2i_1 U1028 ( .x(n3313), .d0(n1978), .sl(n1830), .d1(n1796) );
	mux2i_1 U1029 ( .x(n3314), .d0(n1979), .sl(n1830), .d1(n1797) );
	nand2i_2 U103 ( .x(n1518), .a(n1515), .b(n1519) );
	mux2i_1 U1030 ( .x(n3315), .d0(n1980), .sl(n1830), .d1(n1798) );
	or2_2 U1031 ( .x(n1768), .a(n3935), .b(n3940) );
	mux2_2 U1032 ( .x(n3317), .d0(_RegFile_12__0), .sl(n1829), .d1(WB_data[0]) );
	mux2_2 U1033 ( .x(n3318), .d0(_RegFile_12__1), .sl(n1829), .d1(WB_data[1]) );
	mux2_2 U1034 ( .x(n3319), .d0(_RegFile_12__2), .sl(n1829), .d1(WB_data[2]) );
	mux2_2 U1035 ( .x(n3320), .d0(_RegFile_12__3), .sl(n1829), .d1(WB_data[3]) );
	mux2_2 U1036 ( .x(n3321), .d0(_RegFile_12__4), .sl(n1829), .d1(WB_data[4]) );
	mux2_2 U1037 ( .x(n3322), .d0(_RegFile_12__5), .sl(n1829), .d1(WB_data[5]) );
	mux2_2 U1038 ( .x(n3323), .d0(_RegFile_12__6), .sl(n1829), .d1(WB_data[6]) );
	mux2_2 U1039 ( .x(n3324), .d0(_RegFile_12__7), .sl(n1829), .d1(WB_data[7]) );
	and4i_3 U104 ( .x(n796), .a(n795), .b(___cell__36997_net129977), .c(___cell__36997_net129979),
		.d(___cell__36997_net130187) );
	mux2i_1 U1040 ( .x(n3326), .d0(n1959), .sl(n1829), .d1(n1801) );
	mux2i_1 U1041 ( .x(n3327), .d0(n1936), .sl(n1829), .d1(n1778) );
	mux2i_1 U1042 ( .x(n3328), .d0(n1937), .sl(n1829), .d1(n1779) );
	mux2i_1 U1043 ( .x(n3329), .d0(n1938), .sl(n1829), .d1(n1780) );
	mux2i_1 U1044 ( .x(n3330), .d0(n1939), .sl(n1829), .d1(n1781) );
	mux2i_1 U1045 ( .x(n3331), .d0(n1940), .sl(n1829), .d1(n1782) );
	mux2i_1 U1046 ( .x(n3332), .d0(n1941), .sl(n1829), .d1(n1783) );
	mux2i_1 U1047 ( .x(n3333), .d0(n1942), .sl(n1829), .d1(n1784) );
	mux2i_1 U1048 ( .x(n3334), .d0(n1943), .sl(n1829), .d1(n1785) );
	mux2i_1 U1049 ( .x(n3335), .d0(n1944), .sl(n1829), .d1(n1786) );
	inv_2 U105 ( .x(n694), .a(n693) );
	mux2i_1 U1050 ( .x(n3336), .d0(n1945), .sl(n1829), .d1(n1787) );
	mux2i_1 U1051 ( .x(n3337), .d0(n1946), .sl(n1829), .d1(n1788) );
	mux2i_1 U1052 ( .x(n3338), .d0(n1947), .sl(n1829), .d1(n1789) );
	mux2i_1 U1053 ( .x(n3339), .d0(n1948), .sl(n1829), .d1(n1790) );
	mux2i_1 U1054 ( .x(n3340), .d0(n1949), .sl(n1829), .d1(n1791) );
	mux2i_1 U1055 ( .x(n3341), .d0(n1950), .sl(n1829), .d1(n1792) );
	mux2i_1 U1056 ( .x(n3342), .d0(n1951), .sl(n1829), .d1(n1793) );
	mux2i_1 U1057 ( .x(n3343), .d0(n1952), .sl(n1829), .d1(n1794) );
	mux2i_1 U1058 ( .x(n3344), .d0(n1953), .sl(n1829), .d1(n1795) );
	mux2i_1 U1059 ( .x(n3345), .d0(n1954), .sl(n1829), .d1(n1796) );
	inv_5 U106 ( .x(n704), .a(___cell__36997_net126612) );
	mux2i_1 U1060 ( .x(n3346), .d0(n1955), .sl(n1829), .d1(n1797) );
	buf_3 U1061 ( .x(n959), .a(n957) );
	mux2i_1 U1062 ( .x(n3347), .d0(n1956), .sl(n1829), .d1(n1798) );
	buf_3 U1063 ( .x(n946), .a(n939) );
	or2_2 U1064 ( .x(n1769), .a(n3927), .b(n3940) );
	mux2_2 U1065 ( .x(n3349), .d0(_RegFile_11__0), .sl(n1828), .d1(WB_data[0]) );
	mux2_2 U1066 ( .x(n3350), .d0(_RegFile_11__1), .sl(n1828), .d1(WB_data[1]) );
	mux2_2 U1067 ( .x(n3351), .d0(_RegFile_11__2), .sl(n1828), .d1(WB_data[2]) );
	mux2_2 U1068 ( .x(n3352), .d0(_RegFile_11__3), .sl(n1828), .d1(WB_data[3]) );
	mux2_2 U1069 ( .x(n3353), .d0(_RegFile_11__4), .sl(n1828), .d1(WB_data[4]) );
	nor2i_1 U107 ( .x(n1262), .a(___cell__36997_net126612), .b(n1263) );
	mux2_2 U1070 ( .x(n3354), .d0(_RegFile_11__5), .sl(n1828), .d1(WB_data[5]) );
	mux2_2 U1071 ( .x(n3355), .d0(_RegFile_11__6), .sl(n1828), .d1(WB_data[6]) );
	mux2_2 U1072 ( .x(n3356), .d0(_RegFile_11__7), .sl(n1828), .d1(WB_data[7]) );
	mux2i_1 U1073 ( .x(n3358), .d0(n1935), .sl(n1828), .d1(n1801) );
	mux2i_1 U1074 ( .x(n3359), .d0(n1912), .sl(n1828), .d1(n1778) );
	mux2i_1 U1075 ( .x(n3360), .d0(n1913), .sl(n1828), .d1(n1779) );
	mux2i_1 U1076 ( .x(n3361), .d0(n1914), .sl(n1828), .d1(n1780) );
	mux2i_1 U1077 ( .x(n3362), .d0(n1915), .sl(n1828), .d1(n1781) );
	mux2i_1 U1078 ( .x(n3363), .d0(n1916), .sl(n1828), .d1(n1782) );
	mux2i_1 U1079 ( .x(n3364), .d0(n1917), .sl(n1828), .d1(n1783) );
	oai211_1 U108 ( .x(n1261), .a(n1314), .b(n883), .c(FREEZE), .d(n564) );
	mux2i_1 U1080 ( .x(n3365), .d0(n1918), .sl(n1828), .d1(n1784) );
	mux2i_1 U1081 ( .x(n3366), .d0(n1919), .sl(n1828), .d1(n1785) );
	mux2i_1 U1082 ( .x(n3367), .d0(n1920), .sl(n1828), .d1(n1786) );
	mux2i_1 U1083 ( .x(n3368), .d0(n1921), .sl(n1828), .d1(n1787) );
	mux2i_1 U1084 ( .x(n3369), .d0(n1922), .sl(n1828), .d1(n1788) );
	mux2i_1 U1085 ( .x(n3370), .d0(n1923), .sl(n1828), .d1(n1789) );
	mux2i_1 U1086 ( .x(n3371), .d0(n1924), .sl(n1828), .d1(n1790) );
	mux2i_1 U1087 ( .x(n3372), .d0(n1925), .sl(n1828), .d1(n1791) );
	mux2i_1 U1088 ( .x(n3373), .d0(n1926), .sl(n1828), .d1(n1792) );
	mux2i_1 U1089 ( .x(n3374), .d0(n1927), .sl(n1828), .d1(n1793) );
	nand3_1 U109 ( .x(n3944), .a(WB_index_0), .b(WB_index_4), .c(WB_index_1) );
	mux2i_1 U1090 ( .x(n3375), .d0(n1928), .sl(n1828), .d1(n1794) );
	mux2i_1 U1091 ( .x(n3376), .d0(n1929), .sl(n1828), .d1(n1795) );
	mux2i_1 U1092 ( .x(n3377), .d0(n1930), .sl(n1828), .d1(n1796) );
	mux2i_1 U1093 ( .x(n3378), .d0(n1931), .sl(n1828), .d1(n1797) );
	buf_3 U1094 ( .x(n958), .a(n945) );
	mux2i_1 U1095 ( .x(n3379), .d0(n1932), .sl(n1828), .d1(n1798) );
	or2_2 U1096 ( .x(n1770), .a(n3937), .b(n3939) );
	mux2_2 U1097 ( .x(n3381), .d0(_RegFile_10__0), .sl(n1827), .d1(WB_data[0]) );
	mux2_2 U1098 ( .x(n3382), .d0(_RegFile_10__1), .sl(n1827), .d1(WB_data[1]) );
	mux2_2 U1099 ( .x(n3383), .d0(_RegFile_10__2), .sl(n1827), .d1(WB_data[2]) );
	buf_3 U11 ( .x(reg_out_A[23]), .a(n3958) );
	nand3_1 U110 ( .x(n3943), .a(WB_index_4), .b(n3928), .c(WB_index_1) );
	mux2_2 U1100 ( .x(n3384), .d0(_RegFile_10__3), .sl(n1827), .d1(WB_data[3]) );
	mux2_2 U1101 ( .x(n3385), .d0(_RegFile_10__4), .sl(n1827), .d1(WB_data[4]) );
	mux2_2 U1102 ( .x(n3386), .d0(_RegFile_10__5), .sl(n1827), .d1(WB_data[5]) );
	mux2_2 U1103 ( .x(n3387), .d0(_RegFile_10__6), .sl(n1827), .d1(WB_data[6]) );
	mux2_2 U1104 ( .x(n3388), .d0(_RegFile_10__7), .sl(n1827), .d1(WB_data[7]) );
	mux2i_1 U1105 ( .x(n3390), .d0(n1911), .sl(n1827), .d1(n1801) );
	mux2i_1 U1106 ( .x(n3391), .d0(n1888), .sl(n1827), .d1(n1778) );
	mux2i_1 U1107 ( .x(n3392), .d0(n1889), .sl(n1827), .d1(n1779) );
	mux2i_1 U1108 ( .x(n3393), .d0(n1890), .sl(n1827), .d1(n1780) );
	mux2i_1 U1109 ( .x(n3394), .d0(n1891), .sl(n1827), .d1(n1781) );
	nand3_1 U111 ( .x(n3942), .a(WB_index_4), .b(n3929), .c(WB_index_0) );
	mux2i_1 U1110 ( .x(n3395), .d0(n1892), .sl(n1827), .d1(n1782) );
	mux2i_1 U1111 ( .x(n3396), .d0(n1893), .sl(n1827), .d1(n1783) );
	mux2i_1 U1112 ( .x(n3397), .d0(n1894), .sl(n1827), .d1(n1784) );
	mux2i_1 U1113 ( .x(n3398), .d0(n1895), .sl(n1827), .d1(n1785) );
	mux2i_1 U1114 ( .x(n3399), .d0(n1896), .sl(n1827), .d1(n1786) );
	mux2i_1 U1115 ( .x(n3400), .d0(n1897), .sl(n1827), .d1(n1787) );
	mux2i_1 U1116 ( .x(n3401), .d0(n1898), .sl(n1827), .d1(n1788) );
	mux2i_1 U1117 ( .x(n3402), .d0(n1899), .sl(n1827), .d1(n1789) );
	mux2i_1 U1118 ( .x(n3403), .d0(n1900), .sl(n1827), .d1(n1790) );
	mux2i_1 U1119 ( .x(n3404), .d0(n1901), .sl(n1827), .d1(n1791) );
	nand3_1 U112 ( .x(n3941), .a(n3929), .b(n3928), .c(WB_index_4) );
	mux2i_1 U1120 ( .x(n3405), .d0(n1902), .sl(n1827), .d1(n1792) );
	mux2i_1 U1121 ( .x(n3406), .d0(n1903), .sl(n1827), .d1(n1793) );
	mux2i_1 U1122 ( .x(n3407), .d0(n1904), .sl(n1827), .d1(n1794) );
	mux2i_1 U1123 ( .x(n3408), .d0(n1905), .sl(n1827), .d1(n1795) );
	mux2i_1 U1124 ( .x(n3409), .d0(n1906), .sl(n1827), .d1(n1796) );
	mux2i_1 U1125 ( .x(n3410), .d0(n1907), .sl(n1827), .d1(n1797) );
	mux2i_1 U1126 ( .x(n3411), .d0(n1908), .sl(n1827), .d1(n1798) );
	or2_2 U1127 ( .x(n1771), .a(n3936), .b(n3939) );
	mux2_2 U1128 ( .x(n3413), .d0(_RegFile_9__0), .sl(n1857), .d1(WB_data[0]) );
	mux2_2 U1129 ( .x(n3414), .d0(_RegFile_9__1), .sl(n1857), .d1(WB_data[1]) );
	nand3_1 U113 ( .x(n3940), .a(WB_index_2), .b(WB_index_3), .c(reg_write_WB) );
	mux2_2 U1130 ( .x(n3415), .d0(_RegFile_9__2), .sl(n1857), .d1(WB_data[2]) );
	mux2_2 U1131 ( .x(n3416), .d0(_RegFile_9__3), .sl(n1857), .d1(WB_data[3]) );
	mux2_2 U1132 ( .x(n3417), .d0(_RegFile_9__4), .sl(n1857), .d1(WB_data[4]) );
	mux2_2 U1133 ( .x(n3418), .d0(_RegFile_9__5), .sl(n1857), .d1(WB_data[5]) );
	mux2_2 U1134 ( .x(n3419), .d0(_RegFile_9__6), .sl(n1857), .d1(n691) );
	mux2_2 U1135 ( .x(n3420), .d0(_RegFile_9__7), .sl(n1857), .d1(n692) );
	mux2i_1 U1136 ( .x(n3422), .d0(n2631), .sl(n1857), .d1(n1801) );
	mux2i_1 U1137 ( .x(n3423), .d0(n2608), .sl(n1857), .d1(n1778) );
	mux2i_1 U1138 ( .x(n3424), .d0(n2609), .sl(n1857), .d1(n1779) );
	mux2i_1 U1139 ( .x(n3425), .d0(n2610), .sl(n1857), .d1(n1780) );
	nand3_1 U114 ( .x(n3939), .a(reg_write_WB), .b(n3925), .c(WB_index_3) );
	mux2i_1 U1140 ( .x(n3426), .d0(n2611), .sl(n1857), .d1(n1781) );
	mux2i_1 U1141 ( .x(n3427), .d0(n2612), .sl(n1857), .d1(n1782) );
	mux2i_1 U1142 ( .x(n3428), .d0(n2613), .sl(n1857), .d1(n1783) );
	mux2i_1 U1143 ( .x(n3429), .d0(n2614), .sl(n1857), .d1(n1784) );
	mux2i_1 U1144 ( .x(n3430), .d0(n2615), .sl(n1857), .d1(n1785) );
	mux2i_1 U1145 ( .x(n3431), .d0(n2616), .sl(n1857), .d1(n1786) );
	mux2i_1 U1146 ( .x(n3432), .d0(n2617), .sl(n1857), .d1(n1787) );
	mux2i_1 U1147 ( .x(n3433), .d0(n2618), .sl(n1857), .d1(n1788) );
	mux2i_1 U1148 ( .x(n3434), .d0(n2619), .sl(n1857), .d1(n1789) );
	mux2i_1 U1149 ( .x(n3435), .d0(n2620), .sl(n1857), .d1(n1790) );
	nand3_1 U115 ( .x(n3938), .a(reg_write_WB), .b(n3926), .c(WB_index_2) );
	mux2i_1 U1150 ( .x(n3436), .d0(n2621), .sl(n1857), .d1(n1791) );
	mux2i_1 U1151 ( .x(n3437), .d0(n2622), .sl(n1857), .d1(n1792) );
	mux2i_1 U1152 ( .x(n3438), .d0(n2623), .sl(n1857), .d1(n1793) );
	mux2i_1 U1153 ( .x(n3439), .d0(n2624), .sl(n1857), .d1(n1794) );
	mux2i_1 U1154 ( .x(n3440), .d0(n2625), .sl(n1857), .d1(n1795) );
	mux2i_1 U1155 ( .x(n3441), .d0(n2626), .sl(n1857), .d1(n1796) );
	mux2i_1 U1156 ( .x(n3442), .d0(n2627), .sl(n1857), .d1(n1797) );
	mux2i_1 U1157 ( .x(n3443), .d0(n2628), .sl(n1857), .d1(n1798) );
	or2_2 U1158 ( .x(n1741), .a(n3935), .b(n3939) );
	mux2_2 U1159 ( .x(n3445), .d0(_RegFile_8__0), .sl(n1856), .d1(WB_data[0]) );
	nand3_1 U116 ( .x(n3937), .a(WB_index_0), .b(___cell__6171_net27367), .c(WB_index_1) );
	mux2_2 U1160 ( .x(n3446), .d0(_RegFile_8__1), .sl(n1856), .d1(WB_data[1]) );
	mux2_2 U1161 ( .x(n3447), .d0(_RegFile_8__2), .sl(n1856), .d1(WB_data[2]) );
	mux2_2 U1162 ( .x(n3448), .d0(_RegFile_8__3), .sl(n1856), .d1(WB_data[3]) );
	mux2_2 U1163 ( .x(n3449), .d0(_RegFile_8__4), .sl(n1856), .d1(WB_data[4]) );
	mux2_2 U1164 ( .x(n3450), .d0(_RegFile_8__5), .sl(n1856), .d1(WB_data[5]) );
	mux2_2 U1165 ( .x(n3451), .d0(_RegFile_8__6), .sl(n1856), .d1(n691) );
	mux2_2 U1166 ( .x(n3452), .d0(_RegFile_8__7), .sl(n1856), .d1(WB_data[7]) );
	mux2i_1 U1167 ( .x(n3454), .d0(n2607), .sl(n1856), .d1(n1801) );
	mux2i_1 U1168 ( .x(n3455), .d0(n2584), .sl(n1856), .d1(n1778) );
	mux2i_1 U1169 ( .x(n3456), .d0(n2585), .sl(n1856), .d1(n1779) );
	nand3_1 U117 ( .x(n3936), .a(___cell__6171_net27367), .b(n3928), .c(WB_index_1) );
	mux2i_1 U1170 ( .x(n3457), .d0(n2586), .sl(n1856), .d1(n1780) );
	mux2i_1 U1171 ( .x(n3458), .d0(n2587), .sl(n1856), .d1(n1781) );
	mux2i_1 U1172 ( .x(n3459), .d0(n2588), .sl(n1856), .d1(n1782) );
	mux2i_1 U1173 ( .x(n3460), .d0(n2589), .sl(n1856), .d1(n1783) );
	mux2i_1 U1174 ( .x(n3461), .d0(n2590), .sl(n1856), .d1(n1784) );
	mux2i_1 U1175 ( .x(n3462), .d0(n2591), .sl(n1856), .d1(n1785) );
	mux2i_1 U1176 ( .x(n3463), .d0(n2592), .sl(n1856), .d1(n1786) );
	mux2i_1 U1177 ( .x(n3464), .d0(n2593), .sl(n1856), .d1(n1787) );
	mux2i_1 U1178 ( .x(n3465), .d0(n2594), .sl(n1856), .d1(n1788) );
	mux2i_1 U1179 ( .x(n3466), .d0(n2595), .sl(n1856), .d1(n1789) );
	nand3_1 U118 ( .x(n3935), .a(n3929), .b(___cell__6171_net27367), .c(WB_index_0) );
	mux2i_1 U1180 ( .x(n3467), .d0(n2596), .sl(n1856), .d1(n1790) );
	mux2i_1 U1181 ( .x(n3468), .d0(n2597), .sl(n1856), .d1(n1791) );
	mux2i_1 U1182 ( .x(n3469), .d0(n2598), .sl(n1856), .d1(n1792) );
	mux2i_1 U1183 ( .x(n3470), .d0(n2599), .sl(n1856), .d1(n1793) );
	mux2i_1 U1184 ( .x(n3471), .d0(n2600), .sl(n1856), .d1(n1794) );
	mux2i_1 U1185 ( .x(n3472), .d0(n2601), .sl(n1856), .d1(n1795) );
	mux2i_1 U1186 ( .x(n3473), .d0(n2602), .sl(n1856), .d1(n1796) );
	mux2i_1 U1187 ( .x(n3474), .d0(n2603), .sl(n1856), .d1(n1797) );
	mux2i_1 U1188 ( .x(n3475), .d0(n2604), .sl(n1856), .d1(n1798) );
	buf_3 U1189 ( .x(n920), .a(n989) );
	nand2_2 U119 ( .x(n3934), .a(reg_write_WB), .b(n555) );
	or2_2 U1190 ( .x(n1742), .a(n3927), .b(n3939) );
	mux2_2 U1191 ( .x(n3477), .d0(_RegFile_7__0), .sl(n1855), .d1(WB_data[0]) );
	mux2_2 U1192 ( .x(n3478), .d0(_RegFile_7__1), .sl(n1855), .d1(WB_data[1]) );
	mux2_2 U1193 ( .x(n3479), .d0(_RegFile_7__2), .sl(n1855), .d1(WB_data[2]) );
	mux2_2 U1194 ( .x(n3480), .d0(_RegFile_7__3), .sl(n1855), .d1(WB_data[3]) );
	mux2_2 U1195 ( .x(n3481), .d0(_RegFile_7__4), .sl(n1855), .d1(WB_data[4]) );
	mux2_2 U1196 ( .x(n3482), .d0(_RegFile_7__5), .sl(n1855), .d1(WB_data[5]) );
	mux2_2 U1197 ( .x(n3483), .d0(_RegFile_7__6), .sl(n1855), .d1(WB_data[6]) );
	mux2_2 U1198 ( .x(n3484), .d0(_RegFile_7__7), .sl(n1855), .d1(n692) );
	mux2i_1 U1199 ( .x(n3486), .d0(n2583), .sl(n1855), .d1(n1801) );
	inv_6 U12 ( .x(reg_out_B[12]), .a(n750) );
	nand2i_2 U120 ( .x(n1602), .a(n1395), .b(n1511) );
	mux2i_1 U1200 ( .x(n3487), .d0(n2560), .sl(n1855), .d1(n1778) );
	mux2i_1 U1201 ( .x(n3488), .d0(n2561), .sl(n1855), .d1(n1779) );
	mux2i_1 U1202 ( .x(n3489), .d0(n2562), .sl(n1855), .d1(n1780) );
	mux2i_1 U1203 ( .x(n3490), .d0(n2563), .sl(n1855), .d1(n1781) );
	mux2i_1 U1204 ( .x(n3491), .d0(n2564), .sl(n1855), .d1(n1782) );
	mux2i_1 U1205 ( .x(n3492), .d0(n2565), .sl(n1855), .d1(n1783) );
	mux2i_1 U1206 ( .x(n3493), .d0(n2566), .sl(n1855), .d1(n1784) );
	mux2i_1 U1207 ( .x(n3494), .d0(n2567), .sl(n1855), .d1(n1785) );
	mux2i_1 U1208 ( .x(n3495), .d0(n2568), .sl(n1855), .d1(n1786) );
	mux2i_1 U1209 ( .x(n3496), .d0(n2569), .sl(n1855), .d1(n1787) );
	nand2i_2 U121 ( .x(n1600), .a(n1411), .b(n1511) );
	mux2i_1 U1210 ( .x(n3497), .d0(n2570), .sl(n1855), .d1(n1788) );
	mux2i_1 U1211 ( .x(n3498), .d0(n2571), .sl(n1855), .d1(n1789) );
	mux2i_1 U1212 ( .x(n3499), .d0(n2572), .sl(n1855), .d1(n1790) );
	mux2i_1 U1213 ( .x(n3500), .d0(n2573), .sl(n1855), .d1(n1791) );
	mux2i_1 U1214 ( .x(n3501), .d0(n2574), .sl(n1855), .d1(n1792) );
	mux2i_1 U1215 ( .x(n3502), .d0(n2575), .sl(n1855), .d1(n1793) );
	mux2i_1 U1216 ( .x(n3503), .d0(n2576), .sl(n1855), .d1(n1794) );
	mux2i_1 U1217 ( .x(n3504), .d0(n2577), .sl(n1855), .d1(n1795) );
	mux2i_1 U1218 ( .x(n3505), .d0(n2578), .sl(n1855), .d1(n1796) );
	mux2i_1 U1219 ( .x(n3506), .d0(n2579), .sl(n1855), .d1(n1797) );
	nand2i_2 U122 ( .x(n1648), .a(n1392), .b(n1511) );
	mux2i_1 U1220 ( .x(n3507), .d0(n2580), .sl(n1855), .d1(n1798) );
	or2_2 U1221 ( .x(n1743), .a(n3937), .b(n3938) );
	mux2_2 U1222 ( .x(n3509), .d0(_RegFile_6__0), .sl(n1854), .d1(WB_data[0]) );
	mux2_2 U1223 ( .x(n3510), .d0(_RegFile_6__1), .sl(n1854), .d1(WB_data[1]) );
	mux2_2 U1224 ( .x(n3511), .d0(_RegFile_6__2), .sl(n1854), .d1(WB_data[2]) );
	mux2_2 U1225 ( .x(n3512), .d0(_RegFile_6__3), .sl(n1854), .d1(WB_data[3]) );
	mux2_2 U1226 ( .x(n3513), .d0(_RegFile_6__4), .sl(n1854), .d1(WB_data[4]) );
	mux2_2 U1227 ( .x(n3514), .d0(_RegFile_6__5), .sl(n1854), .d1(WB_data[5]) );
	mux2_2 U1228 ( .x(n3515), .d0(_RegFile_6__6), .sl(n1854), .d1(WB_data[6]) );
	mux2_2 U1229 ( .x(n3516), .d0(_RegFile_6__7), .sl(n1854), .d1(WB_data[7]) );
	nand2i_2 U123 ( .x(n1646), .a(n1354), .b(n1511) );
	mux2i_1 U1230 ( .x(n3518), .d0(n2559), .sl(n1854), .d1(n1801) );
	mux2i_1 U1231 ( .x(n3519), .d0(n2536), .sl(n1854), .d1(n1778) );
	mux2i_1 U1232 ( .x(n3520), .d0(n2537), .sl(n1854), .d1(n1779) );
	mux2i_1 U1233 ( .x(n3521), .d0(n2538), .sl(n1854), .d1(n1780) );
	mux2i_1 U1234 ( .x(n3522), .d0(n2539), .sl(n1854), .d1(n1781) );
	mux2i_1 U1235 ( .x(n3523), .d0(n2540), .sl(n1854), .d1(n1782) );
	mux2i_1 U1236 ( .x(n3524), .d0(n2541), .sl(n1854), .d1(n1783) );
	mux2i_1 U1237 ( .x(n3525), .d0(n2542), .sl(n1854), .d1(n1784) );
	mux2i_1 U1238 ( .x(n3526), .d0(n2543), .sl(n1854), .d1(n1785) );
	mux2i_1 U1239 ( .x(n3527), .d0(n2544), .sl(n1854), .d1(n1786) );
	inv_8 U124 ( .x(n1740), .a(n1511) );
	mux2i_1 U1240 ( .x(n3528), .d0(n2545), .sl(n1854), .d1(n1787) );
	mux2i_1 U1241 ( .x(n3529), .d0(n2546), .sl(n1854), .d1(n1788) );
	mux2i_1 U1242 ( .x(n3530), .d0(n2547), .sl(n1854), .d1(n1789) );
	mux2i_1 U1243 ( .x(n3531), .d0(n2548), .sl(n1854), .d1(n1790) );
	mux2i_1 U1244 ( .x(n3532), .d0(n2549), .sl(n1854), .d1(n1791) );
	mux2i_1 U1245 ( .x(n3533), .d0(n2550), .sl(n1854), .d1(n1792) );
	mux2i_1 U1246 ( .x(n3534), .d0(n2551), .sl(n1854), .d1(n1793) );
	mux2i_1 U1247 ( .x(n3535), .d0(n2552), .sl(n1854), .d1(n1794) );
	mux2i_1 U1248 ( .x(n3536), .d0(n2553), .sl(n1854), .d1(n1795) );
	mux2i_1 U1249 ( .x(n3537), .d0(n2554), .sl(n1854), .d1(n1796) );
	inv_2 U125 ( .x(n1512), .a(n1303) );
	mux2i_1 U1250 ( .x(n3538), .d0(n2555), .sl(n1854), .d1(n1797) );
	mux2i_1 U1251 ( .x(n3539), .d0(n2556), .sl(n1854), .d1(n1798) );
	or2_2 U1252 ( .x(n1744), .a(n3936), .b(n3938) );
	mux2_2 U1253 ( .x(n3541), .d0(_RegFile_5__0), .sl(n1853), .d1(WB_data[0]) );
	mux2_2 U1254 ( .x(n3542), .d0(_RegFile_5__1), .sl(n1853), .d1(WB_data[1]) );
	mux2_2 U1255 ( .x(n3543), .d0(_RegFile_5__2), .sl(n1853), .d1(WB_data[2]) );
	mux2_2 U1256 ( .x(n3544), .d0(_RegFile_5__3), .sl(n1853), .d1(WB_data[3]) );
	mux2_2 U1257 ( .x(n3545), .d0(_RegFile_5__4), .sl(n1853), .d1(WB_data[4]) );
	mux2_2 U1258 ( .x(n3546), .d0(_RegFile_5__5), .sl(n1853), .d1(WB_data[5]) );
	mux2_2 U1259 ( .x(n3547), .d0(_RegFile_5__6), .sl(n1853), .d1(WB_data[6]) );
	nand2i_2 U126 ( .x(n1644), .a(n1400), .b(n1511) );
	mux2_2 U1260 ( .x(n3548), .d0(_RegFile_5__7), .sl(n1853), .d1(WB_data[7]) );
	mux2i_1 U1261 ( .x(n3550), .d0(n2535), .sl(n1853), .d1(n1801) );
	mux2i_1 U1262 ( .x(n3551), .d0(n2512), .sl(n1853), .d1(n1778) );
	mux2i_1 U1263 ( .x(n3552), .d0(n2513), .sl(n1853), .d1(n1779) );
	mux2i_1 U1264 ( .x(n3553), .d0(n2514), .sl(n1853), .d1(n1780) );
	mux2i_1 U1265 ( .x(n3554), .d0(n2515), .sl(n1853), .d1(n1781) );
	mux2i_1 U1266 ( .x(n3555), .d0(n2516), .sl(n1853), .d1(n1782) );
	mux2i_1 U1267 ( .x(n3556), .d0(n2517), .sl(n1853), .d1(n1783) );
	mux2i_1 U1268 ( .x(n3557), .d0(n2518), .sl(n1853), .d1(n1784) );
	mux2i_1 U1269 ( .x(n3558), .d0(n2519), .sl(n1853), .d1(n1785) );
	nand2i_2 U127 ( .x(n1642), .a(n1406), .b(n1511) );
	mux2i_1 U1270 ( .x(n3559), .d0(n2520), .sl(n1853), .d1(n1786) );
	mux2i_1 U1271 ( .x(n3560), .d0(n2521), .sl(n1853), .d1(n1787) );
	mux2i_1 U1272 ( .x(n3561), .d0(n2522), .sl(n1853), .d1(n1788) );
	mux2i_1 U1273 ( .x(n3562), .d0(n2523), .sl(n1853), .d1(n1789) );
	mux2i_1 U1274 ( .x(n3563), .d0(n2524), .sl(n1853), .d1(n1790) );
	mux2i_1 U1275 ( .x(n3564), .d0(n2525), .sl(n1853), .d1(n1791) );
	mux2i_1 U1276 ( .x(n3565), .d0(n2526), .sl(n1853), .d1(n1792) );
	mux2i_1 U1277 ( .x(n3566), .d0(n2527), .sl(n1853), .d1(n1793) );
	mux2i_1 U1278 ( .x(n3567), .d0(n2528), .sl(n1853), .d1(n1794) );
	mux2i_1 U1279 ( .x(n3568), .d0(n2529), .sl(n1853), .d1(n1795) );
	nand2i_2 U128 ( .x(n1640), .a(n1359), .b(n1511) );
	mux2i_1 U1280 ( .x(n3569), .d0(n2530), .sl(n1853), .d1(n1796) );
	mux2i_1 U1281 ( .x(n3570), .d0(n2531), .sl(n1853), .d1(n1797) );
	buf_3 U1282 ( .x(n978), .a(n983) );
	mux2i_1 U1283 ( .x(n3571), .d0(n2532), .sl(n1853), .d1(n1798) );
	or2_2 U1284 ( .x(n1745), .a(n3935), .b(n3938) );
	mux2_2 U1285 ( .x(n3573), .d0(_RegFile_4__0), .sl(n1852), .d1(WB_data[0]) );
	mux2_2 U1286 ( .x(n3574), .d0(_RegFile_4__1), .sl(n1852), .d1(WB_data[1]) );
	mux2_2 U1287 ( .x(n3575), .d0(_RegFile_4__2), .sl(n1852), .d1(WB_data[2]) );
	mux2_2 U1288 ( .x(n3576), .d0(_RegFile_4__3), .sl(n1852), .d1(WB_data[3]) );
	mux2_2 U1289 ( .x(n3577), .d0(_RegFile_4__4), .sl(n1852), .d1(WB_data[4]) );
	nand2i_2 U129 ( .x(n1638), .a(n1304), .b(n1511) );
	mux2_2 U1290 ( .x(n3578), .d0(_RegFile_4__5), .sl(n1852), .d1(WB_data[5]) );
	mux2_2 U1291 ( .x(n3579), .d0(_RegFile_4__6), .sl(n1852), .d1(WB_data[6]) );
	mux2_2 U1292 ( .x(n3580), .d0(_RegFile_4__7), .sl(n1852), .d1(WB_data[7]) );
	buf_3 U1293 ( .x(n924), .a(n937) );
	mux2i_1 U1294 ( .x(n3582), .d0(n2511), .sl(n1852), .d1(n1801) );
	mux2i_1 U1295 ( .x(n3583), .d0(n2488), .sl(n1852), .d1(n1778) );
	mux2i_1 U1296 ( .x(n3584), .d0(n2489), .sl(n1852), .d1(n1779) );
	mux2i_1 U1297 ( .x(n3585), .d0(n2490), .sl(n1852), .d1(n1780) );
	mux2i_1 U1298 ( .x(n3586), .d0(n2491), .sl(n1852), .d1(n1781) );
	mux2i_1 U1299 ( .x(n3587), .d0(n2492), .sl(n1852), .d1(n1782) );
	buf_3 U13 ( .x(Imm[27]), .a(N6382) );
	nand2i_2 U130 ( .x(n1636), .a(n1376), .b(n1303) );
	mux2i_1 U1300 ( .x(n3588), .d0(n2493), .sl(n1852), .d1(n1783) );
	mux2i_1 U1301 ( .x(n3589), .d0(n2494), .sl(n1852), .d1(n1784) );
	mux2i_1 U1302 ( .x(n3590), .d0(n2495), .sl(n1852), .d1(n1785) );
	mux2i_1 U1303 ( .x(n3591), .d0(n2496), .sl(n1852), .d1(n1786) );
	mux2i_1 U1304 ( .x(n3592), .d0(n2497), .sl(n1852), .d1(n1787) );
	mux2i_1 U1305 ( .x(n3593), .d0(n2498), .sl(n1852), .d1(n1788) );
	mux2i_1 U1306 ( .x(n3594), .d0(n2499), .sl(n1852), .d1(n1789) );
	mux2i_1 U1307 ( .x(n3595), .d0(n2500), .sl(n1852), .d1(n1790) );
	mux2i_1 U1308 ( .x(n3596), .d0(n2501), .sl(n1852), .d1(n1791) );
	mux2i_1 U1309 ( .x(n3597), .d0(n2502), .sl(n1852), .d1(n1792) );
	nand2i_2 U131 ( .x(n1634), .a(n1349), .b(n1303) );
	mux2i_1 U1310 ( .x(n3598), .d0(n2503), .sl(n1852), .d1(n1793) );
	mux2i_1 U1311 ( .x(n3599), .d0(n2504), .sl(n1852), .d1(n1794) );
	mux2i_1 U1312 ( .x(n3600), .d0(n2505), .sl(n1852), .d1(n1795) );
	mux2i_1 U1313 ( .x(n3601), .d0(n2506), .sl(n1852), .d1(n1796) );
	mux2i_1 U1314 ( .x(n3602), .d0(n2507), .sl(n1852), .d1(n1797) );
	buf_3 U1315 ( .x(n977), .a(n923) );
	mux2i_1 U1316 ( .x(n3603), .d0(n2508), .sl(n1852), .d1(n1798) );
	buf_3 U1317 ( .x(n925), .a(n937) );
	or2_2 U1318 ( .x(n1746), .a(n3927), .b(n3938) );
	mux2_2 U1319 ( .x(n3605), .d0(_RegFile_3__0), .sl(n1851), .d1(WB_data[0]) );
	nand2i_2 U132 ( .x(n1632), .a(n1340), .b(n1303) );
	buf_3 U1320 ( .x(n927), .a(n936) );
	mux2_2 U1321 ( .x(n3606), .d0(_RegFile_3__1), .sl(n1851), .d1(WB_data[1]) );
	mux2_2 U1322 ( .x(n3607), .d0(_RegFile_3__2), .sl(n1851), .d1(WB_data[2]) );
	mux2_2 U1323 ( .x(n3608), .d0(_RegFile_3__3), .sl(n1851), .d1(WB_data[3]) );
	mux2_2 U1324 ( .x(n3609), .d0(_RegFile_3__4), .sl(n1851), .d1(WB_data[4]) );
	mux2_2 U1325 ( .x(n3610), .d0(_RegFile_3__5), .sl(n1851), .d1(WB_data[5]) );
	mux2_2 U1326 ( .x(n3611), .d0(_RegFile_3__6), .sl(n1851), .d1(WB_data[6]) );
	mux2_2 U1327 ( .x(n3612), .d0(_RegFile_3__7), .sl(n1851), .d1(WB_data[7]) );
	mux2i_1 U1328 ( .x(n3614), .d0(n2487), .sl(n1851), .d1(n1801) );
	mux2i_1 U1329 ( .x(n3615), .d0(n2464), .sl(n1851), .d1(n1778) );
	nand2i_2 U133 ( .x(n1630), .a(n1383), .b(n1303) );
	mux2i_1 U1330 ( .x(n3616), .d0(n2465), .sl(n1851), .d1(n1779) );
	mux2i_1 U1331 ( .x(n3617), .d0(n2466), .sl(n1851), .d1(n1780) );
	mux2i_1 U1332 ( .x(n3618), .d0(n2467), .sl(n1851), .d1(n1781) );
	mux2i_1 U1333 ( .x(n3619), .d0(n2468), .sl(n1851), .d1(n1782) );
	mux2i_1 U1334 ( .x(n3620), .d0(n2469), .sl(n1851), .d1(n1783) );
	mux2i_1 U1335 ( .x(n3621), .d0(n2470), .sl(n1851), .d1(n1784) );
	mux2i_1 U1336 ( .x(n3622), .d0(n2471), .sl(n1851), .d1(n1785) );
	mux2i_1 U1337 ( .x(n3623), .d0(n2472), .sl(n1851), .d1(n1786) );
	mux2i_1 U1338 ( .x(n3624), .d0(n2473), .sl(n1851), .d1(n1787) );
	mux2i_1 U1339 ( .x(n3625), .d0(n2474), .sl(n1851), .d1(n1788) );
	nand2i_2 U134 ( .x(n1628), .a(n1381), .b(n1303) );
	mux2i_1 U1340 ( .x(n3626), .d0(n2475), .sl(n1851), .d1(n1789) );
	mux2i_1 U1341 ( .x(n3627), .d0(n2476), .sl(n1851), .d1(n1790) );
	mux2i_1 U1342 ( .x(n3628), .d0(n2477), .sl(n1851), .d1(n1791) );
	mux2i_1 U1343 ( .x(n3629), .d0(n2478), .sl(n1851), .d1(n1792) );
	mux2i_1 U1344 ( .x(n3630), .d0(n2479), .sl(n1851), .d1(n1793) );
	mux2i_1 U1345 ( .x(n3631), .d0(n2480), .sl(n1851), .d1(n1794) );
	mux2i_1 U1346 ( .x(n3632), .d0(n2481), .sl(n1851), .d1(n1795) );
	mux2i_1 U1347 ( .x(n3633), .d0(n2482), .sl(n1851), .d1(n1796) );
	mux2i_1 U1348 ( .x(n3634), .d0(n2483), .sl(n1851), .d1(n1797) );
	mux2i_1 U1349 ( .x(n3635), .d0(n2484), .sl(n1851), .d1(n1798) );
	nand2i_2 U135 ( .x(n1626), .a(n1379), .b(n1303) );
	or2_2 U1350 ( .x(n1747), .a(n3934), .b(n3937) );
	mux2_2 U1351 ( .x(n3637), .d0(_RegFile_2__0), .sl(n1848), .d1(WB_data[0]) );
	mux2_2 U1352 ( .x(n3638), .d0(_RegFile_2__1), .sl(n1848), .d1(WB_data[1]) );
	mux2_2 U1353 ( .x(n3639), .d0(_RegFile_2__2), .sl(n1848), .d1(WB_data[2]) );
	mux2_2 U1354 ( .x(n3640), .d0(_RegFile_2__3), .sl(n1848), .d1(WB_data[3]) );
	mux2_2 U1355 ( .x(n3641), .d0(_RegFile_2__4), .sl(n1848), .d1(WB_data[4]) );
	mux2_2 U1356 ( .x(n3642), .d0(_RegFile_2__5), .sl(n1848), .d1(WB_data[5]) );
	mux2_2 U1357 ( .x(n3643), .d0(_RegFile_2__6), .sl(n1848), .d1(WB_data[6]) );
	mux2_2 U1358 ( .x(n3644), .d0(_RegFile_2__7), .sl(n1848), .d1(WB_data[7]) );
	mux2i_1 U1359 ( .x(n3646), .d0(n2415), .sl(n1848), .d1(n1801) );
	nand2i_2 U136 ( .x(n1624), .a(n1374), .b(n1303) );
	mux2i_1 U1360 ( .x(n3647), .d0(n2392), .sl(n1848), .d1(n1778) );
	mux2i_1 U1361 ( .x(n3648), .d0(n2393), .sl(n1848), .d1(n1779) );
	mux2i_1 U1362 ( .x(n3649), .d0(n2394), .sl(n1848), .d1(n1780) );
	mux2i_1 U1363 ( .x(n3650), .d0(n2395), .sl(n1848), .d1(n1781) );
	mux2i_1 U1364 ( .x(n3651), .d0(n2396), .sl(n1848), .d1(n1782) );
	buf_3 U1365 ( .x(n930), .a(n987) );
	mux2i_1 U1366 ( .x(n3652), .d0(n2397), .sl(n1848), .d1(n1783) );
	mux2i_1 U1367 ( .x(n3653), .d0(n2398), .sl(n1848), .d1(n1784) );
	mux2i_1 U1368 ( .x(n3654), .d0(n2399), .sl(n1848), .d1(n1785) );
	mux2i_1 U1369 ( .x(n3655), .d0(n2400), .sl(n1848), .d1(n1786) );
	nand2i_2 U137 ( .x(n1622), .a(n1403), .b(n1303) );
	mux2i_1 U1370 ( .x(n3656), .d0(n2401), .sl(n1848), .d1(n1787) );
	mux2i_1 U1371 ( .x(n3657), .d0(n2402), .sl(n1848), .d1(n1788) );
	mux2i_1 U1372 ( .x(n3658), .d0(n2403), .sl(n1848), .d1(n1789) );
	mux2i_1 U1373 ( .x(n3659), .d0(n2404), .sl(n1848), .d1(n1790) );
	mux2i_1 U1374 ( .x(n3660), .d0(n2405), .sl(n1848), .d1(n1791) );
	mux2i_1 U1375 ( .x(n3661), .d0(n2406), .sl(n1848), .d1(n1792) );
	mux2i_1 U1376 ( .x(n3662), .d0(n2407), .sl(n1848), .d1(n1793) );
	mux2i_1 U1377 ( .x(n3663), .d0(n2408), .sl(n1848), .d1(n1794) );
	mux2i_1 U1378 ( .x(n3664), .d0(n2409), .sl(n1848), .d1(n1795) );
	mux2i_1 U1379 ( .x(n3665), .d0(n2410), .sl(n1848), .d1(n1796) );
	nand2i_2 U138 ( .x(n1620), .a(n1409), .b(n1303) );
	mux2i_1 U1380 ( .x(n3666), .d0(n2411), .sl(n1848), .d1(n1797) );
	mux2i_1 U1381 ( .x(n3667), .d0(n2412), .sl(n1848), .d1(n1798) );
	buf_3 U1382 ( .x(n929), .a(n987) );
	or2_2 U1383 ( .x(n1750), .a(n3934), .b(n3936) );
	mux2_2 U1384 ( .x(n3669), .d0(_RegFile_1__0), .sl(n1837), .d1(WB_data[0]) );
	mux2_2 U1385 ( .x(n3670), .d0(_RegFile_1__1), .sl(n1837), .d1(WB_data[1]) );
	mux2_2 U1386 ( .x(n3671), .d0(_RegFile_1__2), .sl(n1837), .d1(WB_data[2]) );
	mux2_2 U1387 ( .x(n3672), .d0(_RegFile_1__3), .sl(n1837), .d1(WB_data[3]) );
	mux2_2 U1388 ( .x(n3673), .d0(_RegFile_1__4), .sl(n1837), .d1(WB_data[4]) );
	mux2_2 U1389 ( .x(n3674), .d0(_RegFile_1__5), .sl(n1837), .d1(WB_data[5]) );
	nand2i_2 U139 ( .x(n1618), .a(n1338), .b(n1303) );
	mux2_2 U1390 ( .x(n3675), .d0(_RegFile_1__6), .sl(n1837), .d1(WB_data[6]) );
	mux2_2 U1391 ( .x(n3676), .d0(_RegFile_1__7), .sl(n1837), .d1(WB_data[7]) );
	inv_2 U1392 ( .x(n1603), .a(n1601) );
	mux2i_1 U1393 ( .x(n3678), .d0(n2151), .sl(n1837), .d1(n1801) );
	mux2i_1 U1394 ( .x(n3679), .d0(n2128), .sl(n1837), .d1(n1778) );
	mux2i_1 U1395 ( .x(n3680), .d0(n2129), .sl(n1837), .d1(n1779) );
	mux2i_1 U1396 ( .x(n3681), .d0(n2130), .sl(n1837), .d1(n1780) );
	mux2i_1 U1397 ( .x(n3682), .d0(n2131), .sl(n1837), .d1(n1781) );
	mux2i_1 U1398 ( .x(n3683), .d0(n2132), .sl(n1837), .d1(n1782) );
	mux2i_1 U1399 ( .x(n3684), .d0(n2133), .sl(n1837), .d1(n1783) );
	exor2_1 U14 ( .x(n3945), .a(n3933), .b(opcode_of_MEM_4) );
	nand2i_2 U140 ( .x(n1616), .a(n1361), .b(n1303) );
	mux2i_1 U1400 ( .x(n3685), .d0(n2134), .sl(n1837), .d1(n1784) );
	mux2i_1 U1401 ( .x(n3686), .d0(n2135), .sl(n1837), .d1(n1785) );
	mux2i_1 U1402 ( .x(n3687), .d0(n2136), .sl(n1837), .d1(n1786) );
	mux2i_1 U1403 ( .x(n3688), .d0(n2137), .sl(n1837), .d1(n1787) );
	mux2i_1 U1404 ( .x(n3689), .d0(n2138), .sl(n1837), .d1(n1788) );
	buf_3 U1405 ( .x(n962), .a(n984) );
	mux2i_1 U1406 ( .x(n3690), .d0(n2139), .sl(n1837), .d1(n1789) );
	mux2i_1 U1407 ( .x(n3691), .d0(n2140), .sl(n1837), .d1(n1790) );
	mux2i_1 U1408 ( .x(n3692), .d0(n2141), .sl(n1837), .d1(n1791) );
	mux2i_1 U1409 ( .x(n3693), .d0(n2142), .sl(n1837), .d1(n1792) );
	nand2i_2 U141 ( .x(n1614), .a(n1346), .b(n1303) );
	mux2i_1 U1410 ( .x(n3694), .d0(n2143), .sl(n1837), .d1(n1793) );
	mux2i_1 U1411 ( .x(n3695), .d0(n2144), .sl(n1837), .d1(n1794) );
	mux2i_1 U1412 ( .x(n3696), .d0(n2145), .sl(n1837), .d1(n1795) );
	mux2i_1 U1413 ( .x(n3697), .d0(n2146), .sl(n1837), .d1(n1796) );
	mux2i_1 U1414 ( .x(n3698), .d0(n2147), .sl(n1837), .d1(n1797) );
	buf_3 U1415 ( .x(n963), .a(n984) );
	mux2i_1 U1416 ( .x(n3699), .d0(n2148), .sl(n1837), .d1(n1798) );
	or2_2 U1417 ( .x(n1761), .a(n3934), .b(n3935) );
	mux2_2 U1418 ( .x(n3701), .d0(_RegFile_0__0), .sl(n1826), .d1(n690) );
	mux2_2 U1419 ( .x(n3702), .d0(_RegFile_0__1), .sl(n1826), .d1(n688) );
	nand2i_2 U142 ( .x(n1612), .a(n1357), .b(n1303) );
	mux2_2 U1420 ( .x(n3703), .d0(_RegFile_0__2), .sl(n1826), .d1(WB_data[2]) );
	mux2_2 U1421 ( .x(n3704), .d0(_RegFile_0__3), .sl(n1826), .d1(WB_data[3]) );
	mux2_2 U1422 ( .x(n3705), .d0(_RegFile_0__4), .sl(n1826), .d1(n687) );
	mux2_2 U1423 ( .x(n3706), .d0(_RegFile_0__5), .sl(n1826), .d1(n689) );
	mux2_2 U1424 ( .x(n3707), .d0(_RegFile_0__6), .sl(n1826), .d1(WB_data[6]) );
	mux2_2 U1425 ( .x(n3708), .d0(_RegFile_0__7), .sl(n1826), .d1(WB_data[7]) );
	inv_2 U1426 ( .x(n1800), .a(n1601) );
	nand2i_2 U1427 ( .x(n1772), .a(n3930), .b(reg_write_WB) );
	mux2i_1 U1428 ( .x(n3733), .d0(n1423), .sl(___cell__36997_net126612), .d1(n1424) );
	mux2i_2 U1429 ( .x(_current_IR_reg_1_net49291), .d0(n800), .sl(___cell__36997_net130681),
		.d1(n801) );
	nand2i_2 U143 ( .x(n1610), .a(n1343), .b(n1303) );
	inv_2 U1430 ( .x(n800), .a(current_IR_1) );
	mux2i_1 U1431 ( .x(n3734), .d0(n1421), .sl(___cell__36997_net126612), .d1(n1422) );
	mux2i_1 U1432 ( .x(n3736), .d0(n1418), .sl(___cell__36997_net126612), .d1(n1419) );
	mux2i_1 U1433 ( .x(n3738), .d0(n631), .sl(___cell__36997_net126612), .d1(n1596) );
	mux2i_1 U1434 ( .x(n3740), .d0(n630), .sl(___cell__36997_net126612), .d1(n1593) );
	mux2i_1 U1435 ( .x(n3741), .d0(n629), .sl(___cell__36997_net130681), .d1(n1592) );
	mux2i_1 U1436 ( .x(n3742), .d0(n632), .sl(___cell__36997_net126612), .d1(n1597) );
	mux2i_1 U1437 ( .x(n3746), .d0(n569), .sl(___cell__36997_net126612), .d1(n1413) );
	mux2i_1 U1438 ( .x(n3748), .d0(n645), .sl(___cell__36997_net126612), .d1(n1330) );
	mux2i_1 U1439 ( .x(n3749), .d0(n1332), .sl(___cell__36997_net130681), .d1(n1333) );
	nand2i_2 U144 ( .x(n1608), .a(n1363), .b(n1303) );
	mux2i_1 U1440 ( .x(n3756), .d0(n1323), .sl(___cell__36997_net130681), .d1(n1324) );
	mux2i_1 U1441 ( .x(n3759), .d0(n1318), .sl(___cell__36997_net126612), .d1(n1319) );
	inv_5 U1442 ( .x(n1319), .a(IR_latched_input[27]) );
	nand2i_2 U1443 ( .x(n1066), .a(n1860), .b(n1718) );
	oai21_1 U1444 ( .x(n3765), .a(n1065), .b(___cell__36997_net126621), .c(n1066) );
	nand2i_2 U1445 ( .x(n1074), .a(n1863), .b(n642) );
	nand2i_2 U1446 ( .x(n1107), .a(n2637), .b(n1718) );
	nand2i_3 U1447 ( .x(n1098), .a(n2635), .b(n1718) );
	nand2i_2 U1448 ( .x(n1086), .a(n2636), .b(n642) );
	oai21_1 U1449 ( .x(n3778), .a(n1065), .b(n1085), .c(n1086) );
	nor3_1 U145 ( .x(n1302), .a(n1303), .b(n1304), .c(n1305) );
	nor2i_1 U1450 ( .x(n1097), .a(n1716), .b(n1485) );
	aoi21_1 U1451 ( .x(n1069), .a(rd_addr[1]), .b(n642), .c(n1719) );
	oai21_1 U1452 ( .x(n3784), .a(n1065), .b(n1061), .c(n1076) );
	aoi21_1 U1453 ( .x(n1076), .a(rd_addr[3]), .b(n642), .c(n1719) );
	aoi21_1 U1454 ( .x(n1070), .a(rd_addr[4]), .b(n1718), .c(n1802) );
	oai21_1 U1455 ( .x(n3785), .a(n1775), .b(n1063), .c(n1070) );
	buf_3 U1456 ( .x(n917), .a(n990) );
	nand2i_2 U1457 ( .x(n1077), .a(n561), .b(n642) );
	nand2i_2 U1458 ( .x(n1122), .a(n671), .b(n1718) );
	inv_5 U1459 ( .x(n1718), .a(n705) );
	nand2i_2 U146 ( .x(n1606), .a(___cell__36997_net129389), .b(n1303) );
	nand2i_2 U1460 ( .x(n1133), .a(n558), .b(n642) );
	oai21_1 U1461 ( .x(n3790), .a(n1132), .b(n1775), .c(n1133) );
	buf_3 U1462 ( .x(n918), .a(n988) );
	buf_3 U1463 ( .x(n919), .a(n988) );
	nand2i_2 U1464 ( .x(n1213), .a(n590), .b(net150785) );
	inv_5 U1465 ( .x(n1650), .a(n1773) );
	inv_2 U1466 ( .x(n856), .a(n340) );
	inv_2 U1467 ( .x(n1682), .a(N504) );
	mux2i_1 U1468 ( .x(n3891), .d0(n1682), .sl(n1650), .d1(___cell__36997_net129389) );
	nor2i_1 U1469 ( .x(n1000), .a(___cell__36997_net130681), .b(n1484) );
	oai21_1 U147 ( .x(n1485), .a(___cell__36997_net127190), .b(n1263), .c(n1307) );
	inv_2 U1470 ( .x(n679), .a(n1000) );
	buf_3 U1471 ( .x(n912), .a(n951) );
	buf_3 U1472 ( .x(n913), .a(n952) );
	inv_2 U1473 ( .x(n1728), .a(reg_dst_of_EX_0) );
	buf_3 U1474 ( .x(n914), .a(n952) );
	inv_2 U1475 ( .x(n801), .a(IR_latched_input[1]) );
	inv_1 U1476 ( .x(n1530), .a(NPC[24]) );
	inv_0 U1477 ( .x(n1529), .a(NPC[25]) );
	and3i_1 U1478 ( .x(PIPEEMPTY), .a(n993), .b(n991), .c(n992) );
	nor2i_1 U1479 ( .x(n991), .a(n1726), .b(n1725) );
	nand2i_2 U148 ( .x(n1716), .a(n2638), .b(n1718) );
	inv_2 U1480 ( .x(n992), .a(n3930) );
	nand2_2 U1481 ( .x(n3930), .a(n3931), .b(n555) );
	inv_2 U1482 ( .x(n3931), .a(n3927) );
	nand2i_2 U1483 ( .x(n993), .a(n1727), .b(n1729) );
	inv_2 U1484 ( .x(n1354), .a(WB_data[11]) );
	inv_2 U1485 ( .x(n1359), .a(WB_data[14]) );
	inv_2 U1486 ( .x(n1383), .a(WB_data[19]) );
	inv_2 U1487 ( .x(n1374), .a(WB_data[22]) );
	inv_2 U1488 ( .x(n1346), .a(WB_data[27]) );
	inv_2 U1489 ( .x(n1343), .a(WB_data[29]) );
	inv_5 U149 ( .x(n843), .a(n847) );
	inv_2 U1490 ( .x(n1532), .a(NPC[22]) );
	inv_2 U1491 ( .x(n1395), .a(WB_data[8]) );
	inv_2 U1492 ( .x(n1552), .a(NPC[1]) );
	inv_2 U1493 ( .x(n1553), .a(NPC[0]) );
	inv_2 U1494 ( .x(n1363), .a(WB_data[30]) );
	inv_2 U1495 ( .x(n1595), .a(IR_latched_input[7]) );
	inv_2 U1496 ( .x(n1594), .a(current_IR_7) );
	inv_2 U1497 ( .x(n1534), .a(NPC[20]) );
	inv_2 U1498 ( .x(n1531), .a(NPC[23]) );
	inv_0 U1499 ( .x(n1536), .a(NPC[18]) );
	buf_14 U15 ( .x(reg_out_A[11]), .a(n3967) );
	inv_2 U150 ( .x(n1316), .a(IR_latched_input[28]) );
	inv_2 U1500 ( .x(n851), .a(IR_latched_input[26]) );
	inv_2 U1501 ( .x(___cell__36997_net129389), .a(WB_data[31]) );
	inv_0 U1502 ( .x(n1535), .a(NPC[19]) );
	inv_2 U1503 ( .x(n1361), .a(WB_data[26]) );
	inv_2 U1504 ( .x(n1439), .a(n4454) );
	inv_1 U1505 ( .x(n1311), .a(Imm[31]) );
	inv_2 U1506 ( .x(n1411), .a(WB_data[9]) );
	inv_2 U1507 ( .x(n1392), .a(WB_data[10]) );
	inv_2 U1508 ( .x(n1400), .a(WB_data[12]) );
	inv_2 U1509 ( .x(n1406), .a(WB_data[13]) );
	and2_3 U151 ( .x(n642), .a(n704), .b(n1461) );
	inv_2 U1510 ( .x(n1304), .a(WB_data[15]) );
	inv_2 U1511 ( .x(n1376), .a(WB_data[16]) );
	inv_2 U1512 ( .x(n1349), .a(WB_data[17]) );
	inv_2 U1513 ( .x(n1340), .a(WB_data[18]) );
	inv_2 U1514 ( .x(n1381), .a(WB_data[20]) );
	inv_2 U1515 ( .x(n1379), .a(WB_data[21]) );
	inv_2 U1516 ( .x(n1403), .a(WB_data[23]) );
	inv_2 U1517 ( .x(n1409), .a(WB_data[24]) );
	inv_2 U1518 ( .x(n1338), .a(WB_data[25]) );
	inv_2 U1519 ( .x(n1357), .a(WB_data[28]) );
	inv_2 U1520 ( .x(n1287), .a(EPC_23) );
	inv_2 U1521 ( .x(n1283), .a(EPC_25) );
	inv_2 U1522 ( .x(n1423), .a(current_IR_0) );
	inv_2 U1523 ( .x(n1421), .a(current_IR_2) );
	inv_5 U1524 ( .x(n1418), .a(current_IR_4) );
	inv_2 U1525 ( .x(n1332), .a(current_IR_17) );
	inv_2 U1526 ( .x(n1323), .a(current_IR_24) );
	inv_5 U1527 ( .x(n1318), .a(current_IR_27) );
	inv_2 U1528 ( .x(n1686), .a(WB_index_1) );
	inv_2 U1529 ( .x(n1424), .a(IR_latched_input[0]) );
	inv_2 U1530 ( .x(n1422), .a(IR_latched_input[2]) );
	inv_2 U1531 ( .x(n1417), .a(IR_latched_input[5]) );
	inv_2 U1532 ( .x(n1596), .a(IR_latched_input[6]) );
	inv_2 U1533 ( .x(n1593), .a(IR_latched_input[8]) );
	inv_2 U1534 ( .x(n1592), .a(IR_latched_input[9]) );
	inv_2 U1535 ( .x(n1416), .a(IR_latched_input[11]) );
	inv_2 U1536 ( .x(n1415), .a(IR_latched_input[12]) );
	inv_2 U1537 ( .x(n1414), .a(IR_latched_input[13]) );
	inv_2 U1538 ( .x(n1413), .a(IR_latched_input[14]) );
	inv_2 U1539 ( .x(n1412), .a(IR_latched_input[15]) );
	inv_2 U1540 ( .x(n1331), .a(IR_latched_input[20]) );
	inv_2 U1541 ( .x(n1324), .a(IR_latched_input[24]) );
	inv_2 U1542 ( .x(n1527), .a(NPC[27]) );
	inv_2 U1543 ( .x(n1526), .a(NPC[28]) );
	inv_2 U1544 ( .x(n1525), .a(NPC[29]) );
	inv_2 U1545 ( .x(n1524), .a(NPC[30]) );
	inv_2 U1546 ( .x(___cell__36997_net129786), .a(NPC[31]) );
	and2_1 U1547 ( .x(n555), .a(n3925), .b(n3926) );
	and2_1 U1548 ( .x(n556), .a(opcode_of_MEM_2), .b(opcode_of_MEM_4) );
	mux2i_1 U1549 ( .x(n628), .d0(n3946), .sl(opcode_of_MEM_1), .d1(n3947) );
	nor2i_6 U155 ( .x(n1691), .a(n772), .b(n340) );
	mux2_6 U1550 ( .x(n637), .d0(n1410), .sl(___cell__36997_net129354), .d1(n1411) );
	mux2_6 U1551 ( .x(n640), .d0(n1380), .sl(___cell__36997_net129354), .d1(n1381) );
	inv_16 U1552 ( .x(n1778), .a(n1647) );
	inv_16 U1553 ( .x(n1779), .a(n1645) );
	inv_16 U1554 ( .x(n1780), .a(n1643) );
	inv_16 U1555 ( .x(n1781), .a(n1641) );
	inv_16 U1556 ( .x(n1782), .a(n1639) );
	inv_16 U1557 ( .x(n1783), .a(n1637) );
	inv_16 U1558 ( .x(n1784), .a(n1635) );
	inv_16 U1559 ( .x(n1785), .a(n1633) );
	inv_5 U156 ( .x(n1071), .a(n339) );
	inv_16 U1560 ( .x(n1786), .a(n1631) );
	inv_16 U1561 ( .x(n1787), .a(n1629) );
	inv_16 U1562 ( .x(n1788), .a(n1627) );
	inv_16 U1563 ( .x(n1789), .a(n1625) );
	inv_16 U1564 ( .x(n1790), .a(n1623) );
	inv_16 U1565 ( .x(n1791), .a(n1621) );
	inv_16 U1566 ( .x(n1792), .a(n1619) );
	inv_16 U1567 ( .x(n1793), .a(n1617) );
	inv_16 U1568 ( .x(n1794), .a(n1615) );
	inv_16 U1569 ( .x(n1795), .a(n1613) );
	and3i_1 U157 ( .x(n1735), .a(n1687), .b(n1575), .c(reg_write_WB) );
	inv_16 U1570 ( .x(n1796), .a(n1611) );
	inv_16 U1571 ( .x(n1797), .a(n1609) );
	inv_16 U1572 ( .x(n1798), .a(n1607) );
	nand2_2 U1573 ( .x(n1604), .a(n1605), .b(n1606) );
	inv_5 U1574 ( .x(n1799), .a(n1604) );
	nand2_2 U1575 ( .x(n1599), .a(n1514), .b(n1600) );
	inv_5 U1576 ( .x(n1801), .a(n1599) );
	inv_16 U1577 ( .x(n1803), .a(n1520) );
	buf_3 U1578 ( .x(n949), .a(n932) );
	buf_3 U1579 ( .x(n950), .a(n932) );
	nand2_2 U158 ( .x(n1734), .a(n1574), .b(n1573) );
	buf_3 U1580 ( .x(n967), .a(n922) );
	buf_3 U1581 ( .x(n966), .a(n922) );
	buf_3 U1582 ( .x(n975), .a(n922) );
	buf_3 U1583 ( .x(n974), .a(n922) );
	buf_3 U1584 ( .x(n976), .a(n923) );
	buf_3 U1585 ( .x(n968), .a(n952) );
	buf_3 U1586 ( .x(n947), .a(n938) );
	buf_3 U1587 ( .x(n969), .a(n952) );
	buf_3 U1588 ( .x(n948), .a(n938) );
	buf_3 U1589 ( .x(n964), .a(n952) );
	exnor2_1 U159 ( .x(n1573), .a(n772), .b(n3926) );
	buf_3 U1590 ( .x(n983), .a(n1858) );
	buf_3 U1591 ( .x(n923), .a(n915) );
	buf_3 U1592 ( .x(n954), .a(n926) );
	buf_3 U1593 ( .x(n972), .a(n986) );
	buf_3 U1594 ( .x(n922), .a(n915) );
	buf_3 U1595 ( .x(n957), .a(n945) );
	buf_3 U1596 ( .x(n945), .a(n939) );
	buf_3 U1597 ( .x(n926), .a(n936) );
	buf_3 U1598 ( .x(n932), .a(n961) );
	buf_3 U1599 ( .x(n938), .a(n961) );
	buf_14 U16 ( .x(Imm[19]), .a(N6366) );
	buf_3 U160 ( .x(n892), .a(n339) );
	buf_3 U1600 ( .x(n939), .a(n961) );
	buf_3 U1601 ( .x(n934), .a(n984) );
	buf_3 U1602 ( .x(n984), .a(n936) );
	buf_3 U1603 ( .x(n961), .a(n988) );
	buf_3 U1604 ( .x(n937), .a(n987) );
	buf_3 U1605 ( .x(n915), .a(n951) );
	buf_3 U1606 ( .x(n988), .a(n921) );
	buf_3 U1607 ( .x(n952), .a(n936) );
	buf_3 U1608 ( .x(n951), .a(n936) );
	buf_3 U1609 ( .x(n987), .a(n921) );
	inv_2 U161 ( .x(n1333), .a(IR_latched_input[17]) );
	buf_3 U1610 ( .x(n970), .a(n972) );
	buf_3 U1611 ( .x(n971), .a(n972) );
	buf_3 U1612 ( .x(n921), .a(n989) );
	buf_3 U1613 ( .x(n990), .a(n970) );
	buf_3 U1614 ( .x(n916), .a(n990) );
	buf_3 U1615 ( .x(n981), .a(n980) );
	buf_3 U1616 ( .x(n989), .a(n971) );
	buf_3 U1617 ( .x(n935), .a(n988) );
	buf_3 U1618 ( .x(n936), .a(n987) );
	buf_3 U1619 ( .x(n980), .a(n983) );
	buf_3 U1620 ( .x(n985), .a(n935) );
	buf_3 U1621 ( .x(n979), .a(n983) );
	buf_3 U1622 ( .x(n982), .a(n964) );
	buf_3 U1623 ( .x(n911), .a(n951) );
	buf_3 U1624 ( .x(n973), .a(n954) );
	buf_3 U1625 ( .x(n953), .a(n926) );
	buf_3 U1626 ( .x(n986), .a(n981) );
	buf_3 U1627 ( .x(n956), .a(n986) );
	buf_3 U1628 ( .x(n955), .a(n986) );
	inv_2 U1631 ( .x(n1330), .a(IR_latched_input[16]) );
	ao22_2 U1633 ( .x(n650), .a(n883), .b(n882), .c(n1517), .d(n881) );
	mux2_5 U1634 ( .x(n653), .d0(n1367), .sl(___cell__36997_net129354), .d1(n1368) );
	inv_2 U1635 ( .x(n335), .a(n879) );
	inv_10 U1637 ( .x(net152024), .a(n728) );
	inv_6 U1638 ( .x(___cell__36997_net130705), .a(net148858) );
	inv_6 U1639 ( .x(net148913), .a(___cell__36997_net130705) );
	inv_2 U1640 ( .x(n1328), .a(IR_latched_input[22]) );
	inv_2 U1641 ( .x(n1326), .a(IR_latched_input[23]) );
	buf_16 U1642 ( .x(reg_out_B[17]), .a(n3978) );
	or2_2 U1644 ( .x(n668), .a(___cell__36997_net129247), .b(n1277) );
	inv_2 U1645 ( .x(n1325), .a(IR_latched_input[21]) );
	inv_12 U1646 ( .x(n1688), .a(n1083) );
	mux2_6 U1647 ( .x(n672), .d0(n1384), .sl(___cell__36997_net129354), .d1(n1385) );
	mux2_6 U1648 ( .x(n673), .d0(n1386), .sl(___cell__36997_net129354), .d1(n1387) );
	mux2_6 U1649 ( .x(n674), .d0(n1339), .sl(___cell__36997_net129354), .d1(n1340) );
	inv_2 U165 ( .x(reg_dst_of_EX_3), .a(n702) );
	mux2i_5 U1650 ( .x(n1336), .d0(n1337), .sl(___cell__36997_net129354), .d1(n1338) );
	inv_7 U1651 ( .x(n698), .a(n1336) );
	nand2_2 U1652 ( .x(n675), .a(___cell__36997_net130713), .b(N6039) );
	inv_2 U1653 ( .x(n693), .a(n333) );
	nand2_2 U1654 ( .x(n676), .a(___cell__36997_net130713), .b(N6040) );
	nand2i_4 U1655 ( .x(n1522), .a(n1523), .b(n1445) );
	inv_7 U1656 ( .x(n744), .a(n1522) );
	nand3i_2 U1657 ( .x(n3948), .a(___cell__36997_net125928), .b(n1000), .c(n744) );
	nand2i_2 U1658 ( .x(n1515), .a(n1516), .b(n1517) );
	or3i_5 U1659 ( .x(n680), .a(n744), .b(___cell__36997_net125928), .c(n679) );
	nand3_1 U166 ( .x(n1727), .a(n1559), .b(n702), .c(n1728) );
	inv_7 U1660 ( .x(___cell__36997_net125928), .a(___cell__36997_net129626) );
	buf_10 U1661 ( .x(reg_out_A[27]), .a(n3954) );
	inv_4 U1662 ( .x(n682), .a(n782) );
	inv_5 U1663 ( .x(n1466), .a(n782) );
	nand4_4 U1664 ( .x(n1706), .a(n639), .b(n640), .c(n1014), .d(n663) );
	nor2_6 U1665 ( .x(n1703), .a(n1701), .b(n1702) );
	nand4_5 U1666 ( .x(n1710), .a(n1128), .b(n637), .c(n1020), .d(n1003) );
	inv_6 U1667 ( .x(n1024), .a(n1344) );
	aoi22_1 U1668 ( .x(n1144), .a(n1344), .b(n797), .c(EPC_27), .d(net150625) );
	inv_0 U1669 ( .x(n683), .a(n847) );
	nand3_1 U167 ( .x(n3927), .a(___cell__6171_net27367), .b(n3928), .c(n3929) );
	inv_6 U1670 ( .x(n847), .a(n850) );
	inv_0 U1671 ( .x(n684), .a(n1377) );
	mux2i_2 U1672 ( .x(n1377), .d0(n1378), .sl(___cell__36997_net129354), .d1(n1379) );
	inv_4 U1673 ( .x(n1014), .a(n1377) );
	inv_2 U1674 ( .x(n685), .a(n1387) );
	inv_2 U1675 ( .x(n1387), .a(WB_data[3]) );
	inv_2 U1676 ( .x(n686), .a(n1390) );
	inv_2 U1677 ( .x(n1390), .a(WB_data[2]) );
	inv_2 U1678 ( .x(n687), .a(n1397) );
	inv_2 U1679 ( .x(n1397), .a(WB_data[4]) );
	nand2i_2 U168 ( .x(n1725), .a(reg_dst_of_MEM_2), .b(n1724) );
	inv_2 U1680 ( .x(n688), .a(n1371) );
	inv_2 U1681 ( .x(n1371), .a(WB_data[1]) );
	inv_2 U1682 ( .x(n689), .a(n1368) );
	inv_2 U1683 ( .x(n1368), .a(WB_data[5]) );
	inv_2 U1684 ( .x(n690), .a(n1366) );
	inv_2 U1685 ( .x(n1366), .a(WB_data[0]) );
	inv_2 U1686 ( .x(n691), .a(n1657) );
	inv_2 U1687 ( .x(n1657), .a(WB_data[6]) );
	inv_2 U1688 ( .x(n692), .a(n1385) );
	inv_2 U1689 ( .x(n1385), .a(WB_data[7]) );
	nor2_1 U169 ( .x(n1724), .a(reg_dst_of_MEM_0), .b(reg_dst_of_MEM_1) );
	buf_14 U1690 ( .x(reg_out_A[28]), .a(n3953) );
	buf_14 U1691 ( .x(reg_out_A[29]), .a(n3952) );
	inv_2 U1693 ( .x(n695), .a(n693) );
	nand2i_2 U1694 ( .x(n1161), .a(n587), .b(net150626) );
	nand2i_2 U1695 ( .x(n1181), .a(n586), .b(net150626) );
	nand2i_2 U1696 ( .x(n1165), .a(n589), .b(net150626) );
	nand2i_2 U1697 ( .x(n1149), .a(n583), .b(net150626) );
	nand2i_2 U1698 ( .x(n1169), .a(n573), .b(net150626) );
	nand2i_2 U1699 ( .x(n1225), .a(n591), .b(net150626) );
	inv_0 U17 ( .x(n1533), .a(NPC[21]) );
	nor2_1 U170 ( .x(n1726), .a(reg_dst_of_MEM_3), .b(reg_dst_of_MEM_4) );
	nand2i_2 U1700 ( .x(n1209), .a(n584), .b(net150626) );
	nand2i_2 U1701 ( .x(n1229), .a(n593), .b(net150626) );
	nand2i_2 U1702 ( .x(n1201), .a(n577), .b(net150626) );
	nand2i_2 U1703 ( .x(n1157), .a(n595), .b(net150626) );
	nand2i_2 U1704 ( .x(n1189), .a(n592), .b(net150626) );
	nand2i_2 U1705 ( .x(n1177), .a(n575), .b(net150626) );
	nand2i_2 U1706 ( .x(n1245), .a(n574), .b(net150626) );
	nand2i_2 U1707 ( .x(n1205), .a(n572), .b(net150626) );
	nand2i_2 U1708 ( .x(n1153), .a(n594), .b(net150626) );
	nand2i_2 U1709 ( .x(n1173), .a(n576), .b(net150626) );
	nand2i_2 U171 ( .x(n1089), .a(n559), .b(n642) );
	inv_5 U1711 ( .x(n1339), .a(N450) );
	inv_10 U1712 ( .x(n697), .a(n1431) );
	nand2i_8 U1713 ( .x(n1431), .a(n1432), .b(n1430) );
	inv_0 U1714 ( .x(n1096), .a(n1431) );
	and2_8 U1715 ( .x(net149679), .a(n780), .b(n787) );
	nand4i_4 U1716 ( .x(n1704), .a(n1372), .b(n1130), .c(n653), .d(n994) );
	nand4_5 U1718 ( .x(n1701), .a(n1024), .b(n1028), .c(n674), .d(n698) );
	inv_0 U1719 ( .x(n699), .a(n1347) );
	nand2i_2 U172 ( .x(n1072), .a(n560), .b(n1718) );
	inv_6 U1720 ( .x(n1009), .a(n1347) );
	mux2i_5 U1721 ( .x(n1347), .d0(n1348), .sl(___cell__36997_net129354), .d1(n1349) );
	nand3_4 U1722 ( .x(n1459), .a(n855), .b(n714), .c(n747) );
	nand4_5 U1723 ( .x(n1702), .a(n1026), .b(n998), .c(n1006), .d(n1009) );
	nand2i_0 U1724 ( .x(n1722), .a(n2634), .b(n1461) );
	nand2i_3 U1725 ( .x(n1143), .a(n1498), .b(n863) );
	nand4i_1 U1727 ( .x(n700), .a(n1456), .b(n1457), .c(n1458), .d(n1444) );
	inv_5 U1728 ( .x(n714), .a(n1455) );
	oai21_1 U1729 ( .x(N6723), .a(n653), .b(n995), .c(n1126) );
	mux2i_1 U173 ( .x(n3737), .d0(n565), .sl(___cell__36997_net130681), .d1(n1417) );
	exnor2_1 U1731 ( .x(___cell__36997_net129977), .a(n1427), .b(n3926) );
	exnor2_1 U1732 ( .x(n1562), .a(n1427), .b(n634) );
	exnor2_2 U1733 ( .x(n1695), .a(n1427), .b(n702) );
	nand2_6 U1734 ( .x(n756), .a(n822), .b(n1446) );
	inv_10 U1736 ( .x(___cell__36997_net125989), .a(___cell__36997_net129381) );
	inv_10 U1737 ( .x(___cell__36997_net125941), .a(___cell__36997_net129378) );
	aoi22_4 U1738 ( .x(n859), .a(n883), .b(n882), .c(n757), .d(n881) );
	inv_6 U1739 ( .x(n757), .a(n752) );
	mux2i_1 U174 ( .x(n3760), .d0(n566), .sl(___cell__36997_net130681), .d1(n1316) );
	exor2_5 U1740 ( .x(n1442), .a(reg_dst_of_EX_4), .b(n1132) );
	exnor2_6 U1741 ( .x(n1570), .a(n1571), .b(n708) );
	mux2i_2 U1743 ( .x(n702), .d0(rd_addr[3]), .sl(n703), .d1(rt_addr[3]) );
	nand2_0 U1744 ( .x(n1731), .a(n3998), .b(n1565) );
	exor2_1 U1745 ( .x(n1685), .a(n1686), .b(n1565) );
	nand2_3 U1747 ( .x(n1432), .a(n739), .b(n815) );
	nand2_8 U1749 ( .x(n705), .a(n704), .b(n1461) );
	mux2i_1 U175 ( .x(n3752), .d0(n567), .sl(___cell__36997_net130681), .d1(n1331) );
	inv_16 U1750 ( .x(n1461), .a(n1260) );
	nand2i_8 U1751 ( .x(n1428), .a(n1315), .b(n1111) );
	inv_0 U1752 ( .x(n707), .a(n683) );
	inv_2 U1753 ( .x(n708), .a(n707) );
	oai21_1 U1754 ( .x(N6718), .a(n3985), .b(___cell__36997_net130580), .c(n996) );
	inv_5 U1755 ( .x(n1337), .a(N443) );
	and2_8 U1756 ( .x(n709), .a(n710), .b(n1694) );
	nor3_2 U1757 ( .x(n710), .a(n333), .b(n715), .c(n761) );
	nand2_1 U1758 ( .x(n1434), .a(n739), .b(n850) );
	nand2_0 U1759 ( .x(n1516), .a(n724), .b(n683) );
	mux2i_1 U176 ( .x(n3747), .d0(n568), .sl(___cell__36997_net130681), .d1(n1412) );
	nand2i_3 U1761 ( .x(n1449), .a(n1446), .b(n822) );
	oai21_1 U1762 ( .x(N6721), .a(n673), .b(n1777), .c(n1238) );
	inv_6 U1763 ( .x(n769), .a(n736) );
	aoi21_1 U1764 ( .x(n1087), .a(rd_addr[2]), .b(n1718), .c(n1802) );
	aoi22_1 U1766 ( .x(n1141), .a(n1355), .b(n797), .c(EPC_28), .d(net150625) );
	mux2i_6 U1767 ( .x(n1355), .d0(n1356), .sl(___cell__36997_net129354), .d1(n1357) );
	nand2i_4 U1768 ( .x(n711), .a(n1429), .b(n753) );
	nand2i_4 U1769 ( .x(n752), .a(n1429), .b(n753) );
	mux2i_1 U177 ( .x(n3745), .d0(n570), .sl(___cell__36997_net130681), .d1(n1414) );
	aoi21_3 U1770 ( .x(n825), .a(n1737), .b(n826), .c(n1451) );
	inv_3 U1771 ( .x(n1500), .a(N5378) );
	aoi21_1 U1772 ( .x(n1075), .a(rd_addr[0]), .b(n1718), .c(n1802) );
	inv_0 U1773 ( .x(n807), .a(n1096) );
	inv_10 U1774 ( .x(n333), .a(n759) );
	mux2i_8 U1775 ( .x(n759), .d0(IR_latched_input[23]), .sl(n760), .d1(current_IR_23) );
	nor2i_2 U1776 ( .x(n1264), .a(n855), .b(n1265) );
	mux2i_8 U1777 ( .x(n712), .d0(n1318), .sl(n728), .d1(n1319) );
	and2_8 U1778 ( .x(n822), .a(n823), .b(n1437) );
	nand2i_0 U1779 ( .x(n713), .a(n1487), .b(n846) );
	mux2i_1 U178 ( .x(n3743), .d0(n571), .sl(___cell__36997_net130681), .d1(n1416) );
	inv_14 U1781 ( .x(n855), .a(n756) );
	nand4i_3 U1782 ( .x(n1455), .a(n1456), .b(n1457), .c(n1458), .d(n1444) );
	nand2_6 U1783 ( .x(___cell__36997_net129632), .a(n812), .b(net148863) );
	oai21_1 U1784 ( .x(N6731), .a(n1003), .b(n995), .c(n1004) );
	inv_8 U1785 ( .x(n1003), .a(n1404) );
	oai21_1 U1786 ( .x(N6719), .a(n1130), .b(n995), .c(n1131) );
	oai211_2 U1789 ( .x(n841), .a(n1081), .b(n843), .c(n767), .d(n724) );
	mux2i_1 U179 ( .x(n2647), .d0(n622), .sl(___cell__36997_net130567), .d1(n845) );
	oai21_1 U1790 ( .x(n3771), .a(n1081), .b(n1775), .c(n1082) );
	nand2i_1 U1791 ( .x(n1491), .a(n1688), .b(n1096) );
	inv_6 U1792 ( .x(n767), .a(n1688) );
	and2_1 U1794 ( .x(n812), .a(n1467), .b(n1688) );
	inv_10 U1795 ( .x(n1437), .a(n1435) );
	inv_2 U1796 ( .x(n717), .a(n1548) );
	inv_0 U1797 ( .x(n718), .a(n715) );
	inv_2 U1798 ( .x(n719), .a(n718) );
	inv_2 U1799 ( .x(n1445), .a(n855) );
	nor2_1 U18 ( .x(n1581), .a(IR_opcode_field[3]), .b(n1321) );
	mux2i_1 U180 ( .x(n2646), .d0(n623), .sl(___cell__36997_net130125), .d1(n871) );
	ao21_4 U1800 ( .x(n721), .a(n1737), .b(n861), .c(n755) );
	exor2_2 U1802 ( .x(n1560), .a(n1561), .b(n759) );
	aoi21_1 U1805 ( .x(n1080), .a(IR_function_field[5]), .b(n1718), .c(n1719) );
	inv_8 U1806 ( .x(n722), .a(N6376) );
	inv_16 U1807 ( .x(Imm[24]), .a(n722) );
	inv_3 U1808 ( .x(n1427), .a(n332) );
	mux2i_2 U181 ( .x(n3763), .d0(n633), .sl(___cell__36997_net130681), .d1(n725) );
	nand2_2 U1810 ( .x(n1137), .a(___cell__36997_net130709), .b(N5449) );
	nand2i_2 U1811 ( .x(n3810), .a(n1101), .b(n1100) );
	nand4_1 U1812 ( .x(n3853), .a(n1139), .b(n668), .c(n1138), .d(n1140) );
	inv_10 U1813 ( .x(n810), .a(NPC[3]) );
	inv_16 U1814 ( .x(n865), .a(NPC[2]) );
	inv_2 U1815 ( .x(n725), .a(n724) );
	inv_2 U1816 ( .x(n726), .a(n1543) );
	oai21_1 U1817 ( .x(N6722), .a(n636), .b(n1777), .c(n1127) );
	oai21_1 U1819 ( .x(N6729), .a(n998), .b(n1777), .c(n999) );
	inv_2 U182 ( .x(n1559), .a(reg_dst_of_EX_4) );
	nor2i_2 U1820 ( .x(n1694), .a(n879), .b(n3990) );
	nand2i_0 U1821 ( .x(n1730), .a(n3998), .b(n3990) );
	oai21_1 U1822 ( .x(n3783), .a(n1774), .b(n1059), .c(n1087) );
	oai21_1 U1823 ( .x(n3766), .a(n1774), .b(n1040), .c(n1079) );
	oai21_1 U1824 ( .x(n3768), .a(n1774), .b(n1043), .c(n1074) );
	oai21_1 U1825 ( .x(n3782), .a(n1774), .b(n1057), .c(n1069) );
	oai21_1 U1826 ( .x(n3786), .a(n856), .b(n1774), .c(n1077) );
	oai21_1 U1827 ( .x(n3789), .a(n772), .b(n1774), .c(n1122) );
	oai21_1 U1828 ( .x(n3773), .a(n3992), .b(n1774), .c(n1112) );
	oai21_1 U1829 ( .x(N6725), .a(n672), .b(n995), .c(n1243) );
	oai21_1 U183 ( .x(n3764), .a(n1065), .b(n1038), .c(n1078) );
	mux2i_8 U1830 ( .x(n1083), .d0(current_IR_30), .sl(net149679), .d1(IR_latched_input[30]) );
	nand2_1 U1831 ( .x(n2707), .a(n729), .b(n1134) );
	inv_2 U1832 ( .x(n729), .a(n742) );
	nor2i_2 U1833 ( .x(n1312), .a(n825), .b(n837) );
	inv_10 U1835 ( .x(n731), .a(n771) );
	inv_10 U1836 ( .x(___cell__36997_net130572), .a(n771) );
	or3i_1 U1837 ( .x(n2706), .a(n1134), .b(n1473), .c(n1090) );
	nand2i_6 U1838 ( .x(n1737), .a(n1689), .b(n1477) );
	nand2i_2 U184 ( .x(n1078), .a(n1859), .b(n642) );
	ao21_3 U1842 ( .x(n733), .a(net150625), .b(EPC_26), .c(n1280) );
	buf_10 U1843 ( .x(net150625), .a(n799) );
	nand2_0 U1844 ( .x(n1110), .a(n1718), .b(IR_opcode_field[5]) );
	mux2i_1 U1845 ( .x(n1479), .d0(n1585), .sl(IR_opcode_field[5]), .d1(n1582) );
	or3i_1 U1846 ( .x(n1438), .a(IR_opcode_field[3]), .b(IR_opcode_field[5]),
		.c(IR_opcode_field[1]) );
	inv_10 U1848 ( .x(n738), .a(n791) );
	inv_10 U1849 ( .x(net148863), .a(n791) );
	mux2i_1 U185 ( .x(n3753), .d0(n646), .sl(___cell__36997_net126612), .d1(n1325) );
	mux2i_8 U1850 ( .x(n739), .d0(IR_latched_input[31]), .sl(net149236), .d1(current_IR_31) );
	nor2_4 U1851 ( .x(n1463), .a(n724), .b(n1578) );
	mux2i_8 U1852 ( .x(n761), .d0(n666), .sl(net149679), .d1(n1327) );
	inv_2 U1853 ( .x(n1327), .a(IR_latched_input[25]) );
	inv_16 U1855 ( .x(net149236), .a(___cell__36997_net130572) );
	nor2i_3 U1856 ( .x(n740), .a(n1590), .b(n741) );
	inv_5 U1857 ( .x(n741), .a(n1454) );
	inv_0 U1858 ( .x(n1591), .a(n1590) );
	oaoi211_1 U1859 ( .x(n742), .a(n745), .b(n744), .c(n743), .d(n883) );
	mux2i_1 U186 ( .x(n3735), .d0(n651), .sl(___cell__36997_net130681), .d1(n1420) );
	inv_2 U1860 ( .x(n743), .a(n1266) );
	inv_0 U1861 ( .x(n745), .a(n1461) );
	nor2i_0 U1862 ( .x(n1266), .a(n1267), .b(___cell__36997_net126612) );
	nand2_5 U1863 ( .x(n835), .a(___cell__36997_net130214), .b(N6023) );
	inv_16 U1864 ( .x(n811), .a(n810) );
	aoi22_2 U1865 ( .x(n1228), .a(N5361), .b(n863), .c(N6028), .d(___cell__36997_net130713) );
	aoi22_2 U1866 ( .x(n1200), .a(N5355), .b(n863), .c(N6022), .d(___cell__36997_net130713) );
	exor2_2 U1867 ( .x(n1696), .a(n1557), .b(n334) );
	inv_10 U1868 ( .x(n1565), .a(n334) );
	mux2i_1 U187 ( .x(n3744), .d0(n652), .sl(___cell__36997_net126612), .d1(n1415) );
	aoi222_1 U1871 ( .x(n1008), .a(NPC[16]), .b(n1802), .c(n1732), .d(EPC_16),
		.e(Cause_Reg_16), .f(n1803) );
	inv_0 U1872 ( .x(n1538), .a(NPC[16]) );
	inv_7 U1873 ( .x(n1736), .a(n1459) );
	nand2i_1 U1875 ( .x(n1483), .a(n1476), .b(n1736) );
	nand2_5 U1876 ( .x(n1489), .a(n1736), .b(n1476) );
	nand4i_5 U1877 ( .x(n1440), .a(n1441), .b(n1444), .c(n1443), .d(n1442) );
	inv_2 U1878 ( .x(n746), .a(n1545) );
	and2_8 U1879 ( .x(n747), .a(n1440), .b(n1313) );
	inv_2 U188 ( .x(n1561), .a(reg_dst_of_EX_2) );
	inv_5 U1881 ( .x(n1517), .a(n711) );
	nor2_3 U1883 ( .x(n1697), .a(n748), .b(n1560) );
	inv_16 U1884 ( .x(n340), .a(n884) );
	inv_10 U1885 ( .x(n1523), .a(n1449) );
	inv_5 U1888 ( .x(n760), .a(net149681) );
	nand2_0 U1889 ( .x(n1084), .a(n642), .b(IR_opcode_field[4]) );
	mux2i_1 U189 ( .x(n3755), .d0(n659), .sl(___cell__36997_net126612), .d1(n1326) );
	nand2_1 U1890 ( .x(n1321), .a(IR_opcode_field[4]), .b(IR_opcode_field[2]) );
	inv_3 U1891 ( .x(n1495), .a(N5382) );
	inv_6 U1892 ( .x(n753), .a(n1428) );
	aoi22_1 U1893 ( .x(n1174), .a(branch_address[5]), .b(n766), .c(N5424),
		.d(___cell__36997_net130709) );
	aoi22_1 U1895 ( .x(n1182), .a(branch_address[17]), .b(n766), .c(N5436),
		.d(___cell__36997_net130709) );
	aoi22_1 U1896 ( .x(n1216), .a(branch_address[15]), .b(n766), .c(N5434),
		.d(___cell__36997_net130709) );
	aoi22_1 U1897 ( .x(n1214), .a(branch_address[13]), .b(n766), .c(N5432),
		.d(___cell__36997_net130709) );
	aoi22_1 U1898 ( .x(n1190), .a(branch_address[11]), .b(n766), .c(N5430),
		.d(___cell__36997_net130709) );
	aoi22_1 U1899 ( .x(n1154), .a(branch_address[1]), .b(n766), .c(N5420),
		.d(___cell__36997_net130709) );
	nor2i_1 U19 ( .x(n1580), .a(n1439), .b(n1568) );
	mux2i_1 U190 ( .x(n3754), .d0(n661), .sl(___cell__36997_net130681), .d1(n1328) );
	aoi21_1 U1900 ( .x(n1178), .a(N5425), .b(___cell__36997_net130709), .c(n1268) );
	or3i_1 U1902 ( .x(n2705), .a(n1134), .b(n1473), .c(n1091) );
	nand2_5 U1903 ( .x(n1446), .a(n1447), .b(___cell__36997_net130306) );
	nand2i_5 U1904 ( .x(n1467), .a(n1468), .b(n1469) );
	inv_1 U1905 ( .x(n1468), .a(n1436) );
	nand4_1 U1906 ( .x(n3852), .a(n1142), .b(n665), .c(n1141), .d(n1143) );
	inv_2 U1907 ( .x(n755), .a(n1479) );
	exnor2_1 U1908 ( .x(n1693), .a(reg_dst_of_EX_2), .b(n338) );
	inv_8 U1909 ( .x(n998), .a(n1352) );
	oai21_1 U191 ( .x(n3769), .a(n1775), .b(n1044), .c(n1080) );
	inv_8 U1910 ( .x(n804), .a(n879) );
	buf_16 U1911 ( .x(Imm[3]), .a(N6334) );
	nand2i_2 U1912 ( .x(n1219), .a(n1006), .b(n797) );
	inv_8 U1913 ( .x(n1006), .a(n1350) );
	mux2i_8 U1915 ( .x(n768), .d0(IR_latched_input[22]), .sl(n769), .d1(n660) );
	nand2i_2 U1916 ( .x(n1183), .a(n699), .b(n797) );
	oai21_1 U1917 ( .x(N6735), .a(n699), .b(n1777), .c(n1010) );
	oai21_1 U1918 ( .x(N6732), .a(___cell__36997_net125941), .b(n1777), .c(n1005) );
	nand2i_2 U1919 ( .x(n1167), .a(___cell__36997_net125941), .b(n797) );
	mux2i_1 U192 ( .x(n3757), .d0(n666), .sl(___cell__36997_net126612), .d1(n1327) );
	oai21_1 U1920 ( .x(N6733), .a(n1006), .b(___cell__36997_net130580), .c(n1007) );
	oai21_1 U1921 ( .x(N6734), .a(n663), .b(n995), .c(n1008) );
	nand2i_2 U1922 ( .x(n1163), .a(n663), .b(n797) );
	mux2i_6 U1923 ( .x(n1341), .d0(n1342), .sl(___cell__36997_net129354), .d1(n1343) );
	nand2i_5 U1924 ( .x(n1106), .a(n1487), .b(n846) );
	nand2i_0 U1925 ( .x(n1085), .a(n1488), .b(n846) );
	inv_10 U1926 ( .x(n846), .a(n841) );
	mux2i_8 U1927 ( .x(n832), .d0(n1418), .sl(n777), .d1(n1419) );
	aoi21_2 U1928 ( .x(n1222), .a(N6036), .b(___cell__36997_net130713), .c(n1295) );
	mux2i_3 U1929 ( .x(n338), .d0(n1334), .sl(net149680), .d1(n1335) );
	mux2i_1 U193 ( .x(n3901), .d0(n1672), .sl(n1650), .d1(n1379) );
	inv_2 U1930 ( .x(n1335), .a(IR_latched_input[18]) );
	aoi22_3 U1931 ( .x(n1212), .a(N5364), .b(n862), .c(N6031), .d(___cell__36997_net130713) );
	inv_16 U1932 ( .x(n862), .a(n1272) );
	exor2_1 U1933 ( .x(n1566), .a(reg_dst_of_MEM_0), .b(n884) );
	exor2_1 U1934 ( .x(n1575), .a(WB_index_0), .b(n856) );
	inv_10 U1935 ( .x(n1477), .a(n1448) );
	nand2_8 U1936 ( .x(n1448), .a(n1106), .b(n1108) );
	mux2i_8 U1937 ( .x(n896), .d0(n1328), .sl(net152024), .d1(n661) );
	inv_2 U1938 ( .x(net152025), .a(net152024) );
	nand2_8 U1939 ( .x(n1429), .a(n716), .b(n1688) );
	inv_2 U194 ( .x(n1672), .a(N514) );
	nand2i_4 U1940 ( .x(n1236), .a(n1508), .b(n862) );
	inv_16 U1941 ( .x(n797), .a(___cell__36997_net129632) );
	or2_3 U1943 ( .x(n758), .a(net151343), .b(n662) );
	inv_0 U1944 ( .x(net151343), .a(n799) );
	and2_6 U1945 ( .x(n867), .a(n868), .b(net148863) );
	mux2i_5 U1946 ( .x(n772), .d0(IR_latched_input[19]), .sl(n760), .d1(current_IR_19) );
	inv_2 U1947 ( .x(n1016), .a(n1372) );
	or2_4 U1948 ( .x(n1100), .a(n1733), .b(n1037) );
	or2_8 U1949 ( .x(n764), .a(n1733), .b(n1037) );
	mux2i_1 U195 ( .x(n3922), .d0(n1649), .sl(n1650), .d1(n1366) );
	or2_8 U1950 ( .x(n763), .a(n1733), .b(n1037) );
	nand2i_2 U1951 ( .x(n1733), .a(n1309), .b(n887) );
	oai21_5 U1952 ( .x(n1037), .a(n1484), .b(n1480), .c(n1554) );
	inv_3 U1953 ( .x(n1497), .a(N6047) );
	oai21_1 U1955 ( .x(n1804), .a(___cell__36997_net129624), .b(___cell__36997_net129625),
		.c(___cell__36997_net130681) );
	mux2i_8 U1956 ( .x(n332), .d0(n1324), .sl(net149236), .d1(n1323) );
	oai21_1 U1957 ( .x(n3777), .a(n1094), .b(n1085), .c(n1098) );
	nand2i_2 U1958 ( .x(n1094), .a(___cell__36997_net127190), .b(n1480) );
	oai21_1 U1959 ( .x(n3772), .a(n1113), .b(n1065), .c(n1114) );
	inv_2 U196 ( .x(n1649), .a(N535) );
	oai21_1 U1960 ( .x(n1488), .a(n1081), .b(n1113), .c(n3992) );
	aoi22_2 U1961 ( .x(n1152), .a(N5352), .b(n895), .c(N6019), .d(___cell__36997_net130214) );
	mux2i_8 U1964 ( .x(IR_latched_1), .d0(n801), .sl(net149236), .d1(n800) );
	buf_10 U1965 ( .x(reg_out_A[22]), .a(n3959) );
	ao22_6 U1968 ( .x(___cell__36997_net129524), .a(n721), .b(n1523), .c(n855),
		.d(n740) );
	mux2i_1 U197 ( .x(n3911), .d0(n1662), .sl(n1650), .d1(n1354) );
	or2_8 U1970 ( .x(n771), .a(n3949), .b(n3950) );
	mux2i_1 U1971 ( .x(n3750), .d0(n1334), .sl(___cell__36997_net126612), .d1(n1335) );
	inv_2 U1972 ( .x(n1334), .a(current_IR_18) );
	inv_10 U1973 ( .x(n337), .a(n772) );
	inv_0 U1974 ( .x(n1329), .a(IR_latched_input[19]) );
	buf_16 U1975 ( .x(reg_out_A[9]), .a(n3969) );
	oai21_1 U1976 ( .x(n773), .a(n1317), .b(n847), .c(n1688) );
	inv_0 U1978 ( .x(n842), .a(n1688) );
	inv_2 U198 ( .x(n1662), .a(N524) );
	inv_4 U1980 ( .x(counter[1]), .a(n780) );
	oai21_4 U1981 ( .x(n1065), .a(n1484), .b(n1480), .c(___cell__36997_net130681) );
	oai21_4 U1982 ( .x(n1775), .a(n1484), .b(n1480), .c(___cell__36997_net126612) );
	oai21_4 U1983 ( .x(n1774), .a(n1484), .b(n1480), .c(___cell__36997_net130681) );
	oai21_2 U1984 ( .x(n854), .a(n1484), .b(n1480), .c(n1554) );
	nor2i_0 U1985 ( .x(n1268), .a(branch_address[6]), .b(n738) );
	oai21_1 U1986 ( .x(n1237), .a(n738), .b(n1722), .c(___cell__36997_net126604) );
	nor2i_0 U1987 ( .x(n1278), .a(branch_address[29]), .b(n738) );
	mux2i_1 U1988 ( .x(n1598), .d0(n2633), .sl(n738), .d1(n1471) );
	nor2i_0 U1989 ( .x(n1280), .a(branch_address[26]), .b(n738) );
	inv_2 U199 ( .x(n1499), .a(N5446) );
	inv_0 U1991 ( .x(n776), .a(net149680) );
	inv_2 U1992 ( .x(n777), .a(n776) );
	aoi22_2 U1993 ( .x(n1147), .a(branch_address[27]), .b(n766), .c(N6045),
		.d(___cell__36997_net130713) );
	inv_14 U1994 ( .x(___cell__36997_net130713), .a(___cell__36997_net129239) );
	nor2i_1 U1995 ( .x(n1300), .a(N6029), .b(___cell__36997_net129239) );
	inv_2 U1997 ( .x(n783), .a(___cell__36997_net129247) );
	nand4_1 U1998 ( .x(n3842), .a(n1222), .b(n784), .c(n1223), .d(n1221) );
	inv_5 U1999 ( .x(n784), .a(n1220) );
	inv_4 U20 ( .x(n1067), .a(n850) );
	mux2i_1 U200 ( .x(n3902), .d0(n1671), .sl(n1650), .d1(n1381) );
	nand2i_4 U2000 ( .x(n1490), .a(n785), .b(n1699) );
	inv_3 U2001 ( .x(n785), .a(n855) );
	exnor2_3 U2002 ( .x(n1684), .a(n655), .b(n333) );
	mux2i_3 U2003 ( .x(n818), .d0(n773), .sl(n1578), .d1(n3989) );
	aoi222_1 U2004 ( .x(n1007), .a(NPC[15]), .b(n1719), .c(n1732), .d(EPC_15),
		.e(Cause_Reg_15), .f(n1803) );
	inv_0 U2005 ( .x(n1539), .a(NPC[15]) );
	oaoi211_1 U2006 ( .x(_counter_reg_0_net48671), .a(___cell__36997_net127189),
		.b(___cell__36997_net127190), .c(n777), .d(counter[0]) );
	nor2i_0 U2007 ( .x(_counter_reg_1_net48651), .a(n790), .b(n4011) );
	buf_1 U2008 ( .x(n790), .a(counter[1]) );
	nand2i_8 U2009 ( .x(___cell__36997_net129247), .a(___cell__36997_net129626),
		.b(n738) );
	inv_2 U201 ( .x(n1671), .a(N515) );
	oai21_6 U2010 ( .x(n791), .a(___cell__36997_net129624), .b(___cell__36997_net129625),
		.c(___cell__36997_net130681) );
	inv_16 U2011 ( .x(___cell__36997_net130681), .a(___cell__36997_net127190) );
	inv_10 U2012 ( .x(___cell__36997_net130214), .a(___cell__36997_net129239) );
	buf_16 U2014 ( .x(net150626), .a(n799) );
	inv_16 U2015 ( .x(___cell__36997_net129354), .a(n798) );
	exor2_3 U2017 ( .x(n795), .a(___cell__6171_net27367), .b(___cell__36997_net129477) );
	inv_0 U2018 ( .x(___cell__36997_net126621), .a(IR_latched_1) );
	inv_10 U2019 ( .x(n1578), .a(n1111) );
	nor2i_1 U202 ( .x(n1109), .a(n1717), .b(n1485) );
	buf_16 U2020 ( .x(n802), .a(n1258) );
	oai21_1 U2021 ( .x(n3774), .a(n842), .b(n1775), .c(n1084) );
	mux2i_1 U2022 ( .x(n3762), .d0(n658), .sl(___cell__36997_net126612), .d1(n842) );
	and4i_1 U2023 ( .x(n1309), .a(n1310), .b(n842), .c(n725), .d(n683) );
	nand2_6 U2024 ( .x(n1435), .a(n859), .b(n1436) );
	buf_16 U2026 ( .x(reg_out_A[26]), .a(n3955) );
	buf_14 U2027 ( .x(n878), .a(n889) );
	inv_2 U2028 ( .x(n808), .a(n807) );
	inv_2 U2029 ( .x(n1496), .a(N6048) );
	oai21_1 U203 ( .x(n3780), .a(n1775), .b(n1108), .c(n1109) );
	inv_7 U2030 ( .x(n809), .a(n1051) );
	inv_10 U2031 ( .x(IR_latched_8), .a(n1049) );
	aoi222_1 U2032 ( .x(n1010), .a(NPC[17]), .b(n1719), .c(n1732), .d(EPC_17),
		.e(Cause_Reg_17), .f(n1803) );
	inv_0 U2033 ( .x(n1537), .a(NPC[17]) );
	nand2_8 U2035 ( .x(___cell__36997_net127155), .a(net148863), .b(n1492) );
	aoi22_1 U2036 ( .x(n1240), .a(branch_address[3]), .b(n766), .c(N6021),
		.d(___cell__36997_net130713) );
	nand2i_2 U2037 ( .x(n1140), .a(n1497), .b(___cell__36997_net130713) );
	nand2i_2 U2038 ( .x(n1198), .a(n1505), .b(___cell__36997_net130713) );
	nand2i_2 U2039 ( .x(n1217), .a(n1510), .b(___cell__36997_net130713) );
	oai21_1 U204 ( .x(n3767), .a(n1065), .b(n1041), .c(n1073) );
	aoi22_1 U2040 ( .x(n1255), .a(branch_address[2]), .b(net148865), .c(N6020),
		.d(___cell__36997_net130713) );
	nand2i_2 U2041 ( .x(n1250), .a(n1501), .b(___cell__36997_net130713) );
	nand2i_2 U2043 ( .x(n1194), .a(n1507), .b(___cell__36997_net130713) );
	nand2i_2 U2044 ( .x(n1136), .a(n1496), .b(___cell__36997_net130713) );
	nor2_3 U2046 ( .x(n1293), .a(net148916), .b(n1294) );
	nor2_3 U2047 ( .x(n1275), .a(net148916), .b(n1276) );
	nor2_4 U2048 ( .x(n1282), .a(net148916), .b(n1283) );
	inv_3 U2049 ( .x(net150785), .a(net148916) );
	nand2i_2 U205 ( .x(n1073), .a(n1862), .b(n1718) );
	inv_14 U2050 ( .x(net148916), .a(___cell__36997_net130217) );
	mux2i_1 U2051 ( .x(n849), .d0(current_IR_3), .sl(n731), .d1(IR_latched_input[3]) );
	inv_0 U2052 ( .x(n1546), .a(NPC[8]) );
	aoi222_1 U2053 ( .x(n1032), .a(NPC[8]), .b(n1802), .c(n1732), .d(EPC_8),
		.e(Cause_Reg_8), .f(n1803) );
	inv_0 U2054 ( .x(n1551), .a(n866) );
	aoi222_1 U2055 ( .x(n1253), .a(n737), .b(n1719), .c(n1732), .d(EPC_2),
		.e(Cause_Reg_2), .f(n1803) );
	mux2i_1 U2056 ( .x(n1091), .d0(n1588), .sl(slot_num_0), .d1(n1589) );
	exnor2_1 U2057 ( .x(n1314), .a(slot_num_1), .b(slot_num_0) );
	nand2i_0 U2058 ( .x(n1267), .a(slot_num_1), .b(slot_num_0) );
	nand2_2 U2059 ( .x(n1576), .a(slot_num_1), .b(slot_num_0) );
	inv_2 U206 ( .x(n1059), .a(IR_latched_13) );
	nor2i_1 U2060 ( .x(n1714), .a(slot_num_0), .b(n557) );
	buf_16 U2061 ( .x(reg_out_A[5]), .a(n3972) );
	inv_0 U2062 ( .x(n1047), .a(n817) );
	inv_0 U2064 ( .x(n820), .a(n809) );
	buf_16 U2065 ( .x(Imm[7]), .a(N6342) );
	inv_2 U2066 ( .x(n861), .a(n1438) );
	mux2i_1 U2067 ( .x(n3758), .d0(n852), .sl(___cell__36997_net130681), .d1(n1067) );
	oai21_1 U2068 ( .x(n3770), .a(n1067), .b(n1774), .c(n1068) );
	inv_5 U2069 ( .x(n1426), .a(n333) );
	oai21_1 U207 ( .x(n3781), .a(n1775), .b(n1055), .c(n1075) );
	nor2_0 U2070 ( .x(n1519), .a(n1730), .b(n1425) );
	nor2_0 U2071 ( .x(n1521), .a(n1731), .b(n1425) );
	nand2i_0 U2072 ( .x(n1712), .a(___cell__36997_net125928), .b(n1713) );
	inv_10 U2073 ( .x(n1713), .a(n1467) );
	inv_2 U2074 ( .x(n826), .a(n1474) );
	inv_5 U2075 ( .x(n1475), .a(n1451) );
	nand2i_2 U2076 ( .x(n1474), .a(opcode_of_MEM_1), .b(n1690) );
	nand2_1 U2077 ( .x(n1487), .a(n1578), .b(n1113) );
	nand2_0 U2078 ( .x(n1310), .a(n1578), .b(n1113) );
	nand3_0 U2079 ( .x(n1425), .a(n1426), .b(n1427), .c(___cell__36997_net129477) );
	nand2i_2 U208 ( .x(n1039), .a(n720), .b(n1718) );
	ao21_1 U2081 ( .x(n2708), .a(___cell__36997_net130681), .b(n1035), .c(n1036) );
	and3i_5 U2082 ( .x(n834), .a(net151366), .b(n1489), .c(n1490) );
	inv_0 U2083 ( .x(n1035), .a(n834) );
	inv_10 U2084 ( .x(net151366), .a(___cell__36997_net127189) );
	inv_10 U2085 ( .x(___cell__36997_net127189), .a(___cell__36997_net129524) );
	inv_0 U2087 ( .x(n836), .a(n840) );
	inv_3 U2088 ( .x(n840), .a(n1462) );
	mux2i_6 U2089 ( .x(reg_dst_of_EX_2), .d0(n559), .sl(reg_dst), .d1(n670) );
	nor2_1 U209 ( .x(n1104), .a(n1776), .b(n654) );
	inv_0 U2090 ( .x(n1044), .a(n888) );
	inv_0 U2091 ( .x(n1308), .a(NPC[6]) );
	oai21_1 U2092 ( .x(n3776), .a(n1094), .b(n713), .c(n1107) );
	inv_0 U2093 ( .x(n1095), .a(n713) );
	buf_16 U2094 ( .x(Imm[21]), .a(N6370) );
	ao221_4 U2095 ( .x(n1689), .a(n1430), .b(n846), .c(n818), .d(n739), .e(n840) );
	nand3i_3 U2096 ( .x(n1462), .a(n712), .b(n1463), .c(n1464) );
	inv_10 U2097 ( .x(n1430), .a(n1428) );
	mux2i_8 U2098 ( .x(n1317), .d0(n1318), .sl(n728), .d1(n1319) );
	exor2_2 U2099 ( .x(n1567), .a(n1088), .b(reg_dst_of_MEM_2) );
	buf_14 U21 ( .x(Imm[9]), .a(N6346) );
	nand2i_2 U210 ( .x(n3815), .a(n1104), .b(n763) );
	exor2_1 U2100 ( .x(n1574), .a(WB_index_2), .b(n1088) );
	oai21_1 U2101 ( .x(n3788), .a(n3986), .b(n1065), .c(n1089) );
	nand4_5 U2102 ( .x(n1444), .a(n1088), .b(n1071), .c(n1691), .d(n1132) );
	buf_14 U2104 ( .x(n888), .a(IR_latched_5) );
	aoi22_1 U2105 ( .x(n1138), .a(n1341), .b(n797), .c(EPC_29), .d(net150625) );
	aoi222_1 U2106 ( .x(n1004), .a(NPC[13]), .b(n1719), .c(n1732), .d(EPC_13),
		.e(Cause_Reg_13), .f(n1803) );
	inv_0 U2107 ( .x(n1541), .a(NPC[13]) );
	oai31_1 U2108 ( .x(n3779), .a(n1094), .b(n1095), .c(n808), .d(n1097) );
	nand2_6 U2109 ( .x(n1469), .a(n1466), .b(n808) );
	mux2i_1 U211 ( .x(n3892), .d0(n1681), .sl(n1650), .d1(n1363) );
	nand2i_8 U2110 ( .x(n1436), .a(n1067), .b(n697) );
	aoi222_1 U2111 ( .x(n1011), .a(NPC[18]), .b(n1802), .c(n1732), .d(EPC_18),
		.e(Cause_Reg_18), .f(n1803) );
	inv_0 U2112 ( .x(n1055), .a(IR_latched_11) );
	aoi21_2 U2113 ( .x(n1172), .a(N5356), .b(n862), .c(n1270) );
	nand4_1 U2114 ( .x(n3847), .a(n1193), .b(n1192), .c(n1194), .d(n1195) );
	nand4_3 U2115 ( .x(n1571), .a(n1711), .b(n1708), .c(n1705), .d(n1703) );
	buf_16 U2116 ( .x(Imm[26]), .a(N6380) );
	aoi22_2 U2117 ( .x(n1218), .a(N5366), .b(n895), .c(EPC_15), .d(net150625) );
	buf_16 U2118 ( .x(reg_out_A[10]), .a(n3968) );
	nand3i_1 U2119 ( .x(n3823), .a(n1237), .b(net148916), .c(n1134) );
	inv_2 U212 ( .x(n1681), .a(N505) );
	mux2i_8 U2120 ( .x(n850), .d0(n851), .sl(net149236), .d1(n852) );
	nand4i_2 U2121 ( .x(n3827), .a(n1239), .b(n1240), .c(n1241), .d(n1242) );
	nand4i_2 U2122 ( .x(n3826), .a(n1254), .b(n1255), .c(n1256), .d(n1257) );
	mux2i_8 U2123 ( .x(IR_latched_12), .d0(n1415), .sl(net149236), .d1(n652) );
	nor2_4 U2125 ( .x(n1284), .a(net148913), .b(n1285) );
	inv_0 U2126 ( .x(n1549), .a(NPC[4]) );
	aoi222_1 U2127 ( .x(n1127), .a(NPC[4]), .b(n1719), .c(n1732), .d(EPC_4),
		.e(Cause_Reg_4), .f(n1803) );
	aoi222_1 U2128 ( .x(n1005), .a(NPC[14]), .b(n1802), .c(n1732), .d(EPC_14),
		.e(Cause_Reg_14), .f(n1803) );
	inv_0 U2129 ( .x(n1540), .a(NPC[14]) );
	or2_4 U213 ( .x(n665), .a(___cell__36997_net129247), .b(n1279) );
	aoi222_1 U2130 ( .x(n1238), .a(n811), .b(n1802), .c(n1732), .d(EPC_3),
		.e(Cause_Reg_3), .f(n1803) );
	inv_0 U2131 ( .x(n1550), .a(n811) );
	nand2i_2 U2132 ( .x(n1482), .a(n721), .b(n1523) );
	mux2i_2 U2133 ( .x(n1315), .d0(n566), .sl(n731), .d1(n1316) );
	inv_5 U2134 ( .x(n857), .a(n856) );
	inv_0 U2135 ( .x(n1544), .a(NPC[10]) );
	aoi222_1 U2136 ( .x(n997), .a(NPC[10]), .b(n1802), .c(n1732), .d(EPC_10),
		.e(Cause_Reg_10), .f(n1803) );
	nand2i_1 U2137 ( .x(n1192), .a(n1018), .b(n797) );
	nand2i_1 U2138 ( .x(n1196), .a(n1020), .b(n797) );
	nand2i_1 U2139 ( .x(n1235), .a(n1016), .b(n797) );
	inv_2 U214 ( .x(n1279), .a(N5447) );
	nand2i_1 U2140 ( .x(n1150), .a(n640), .b(n797) );
	nand2i_1 U2141 ( .x(n1233), .a(n1014), .b(n797) );
	nand2i_1 U2142 ( .x(n1191), .a(n998), .b(n797) );
	nand2i_1 U2143 ( .x(n1159), .a(n3985), .b(n797) );
	nand2i_1 U2144 ( .x(n1247), .a(n672), .b(n797) );
	nand2i_1 U2145 ( .x(n1175), .a(n653), .b(n797) );
	nand2i_1 U2146 ( .x(n1179), .a(n1128), .b(n797) );
	nand2i_2 U2147 ( .x(n1257), .a(n1252), .b(n797) );
	nand2i_2 U2148 ( .x(n1242), .a(n673), .b(n797) );
	nand2i_2 U2149 ( .x(n1223), .a(n674), .b(n797) );
	mux2i_1 U215 ( .x(n3913), .d0(n1660), .sl(n1650), .d1(n1411) );
	nand2i_1 U2150 ( .x(n1203), .a(n636), .b(n797) );
	nand2i_1 U2151 ( .x(n1171), .a(n1031), .b(n797) );
	nand2i_1 U2152 ( .x(n1215), .a(n1003), .b(n797) );
	nand2i_1 U2153 ( .x(n1231), .a(n638), .b(n797) );
	nand2i_1 U2154 ( .x(n1211), .a(n639), .b(n797) );
	nand2i_1 U2155 ( .x(n1155), .a(n1130), .b(n797) );
	nand2i_1 U2156 ( .x(n1227), .a(n1001), .b(n797) );
	nand2i_1 U2157 ( .x(n1207), .a(n637), .b(n797) );
	aoi22_1 U2158 ( .x(n1248), .a(___cell__36997_net129381), .b(n797), .c(N5445),
		.d(___cell__36997_net130709) );
	buf_16 U2159 ( .x(reg_out_A[25]), .a(n3956) );
	inv_2 U216 ( .x(n1660), .a(N526) );
	aoi22_1 U2160 ( .x(n860), .a(n883), .b(n882), .c(n1517), .d(n881) );
	nand4_1 U2161 ( .x(n3845), .a(n1232), .b(n675), .c(n1233), .d(n1234) );
	oai22_1 U2162 ( .x(n3791), .a(n705), .b(n813), .c(n854), .d(n1038) );
	oai21_1 U2163 ( .x(n3792), .a(n3995), .b(___cell__36997_net126621), .c(n1039) );
	oai22_1 U2164 ( .x(n3793), .a(n1776), .b(n870), .c(n3995), .d(n1040) );
	oai21_1 U2165 ( .x(n3794), .a(n3995), .b(n1041), .c(n1042) );
	oai22_1 U2167 ( .x(n3796), .a(n1776), .b(n845), .c(n3995), .d(n1044) );
	oai21_1 U2168 ( .x(n3797), .a(n1045), .b(n3995), .c(n1046) );
	oai21_1 U2169 ( .x(n3798), .a(n1047), .b(n3995), .c(n1048) );
	inv_2 U217 ( .x(n1680), .a(N506) );
	oai21_1 U2170 ( .x(n3799), .a(n1049), .b(n3995), .c(n1050) );
	oai21_1 U2171 ( .x(n3800), .a(n820), .b(n3995), .c(n1052) );
	oai21_1 U2172 ( .x(n3803), .a(n1057), .b(n854), .c(n1058) );
	oai21_1 U2173 ( .x(n3804), .a(n1059), .b(n854), .c(n1060) );
	oai21_1 U2174 ( .x(n3806), .a(n1063), .b(n3995), .c(n1064) );
	oai21_1 U2175 ( .x(n3805), .a(n1061), .b(n854), .c(n1062) );
	inv_16 U2176 ( .x(n863), .a(n1272) );
	inv_16 U2177 ( .x(n1272), .a(n867) );
	mux2i_8 U2178 ( .x(IR_latched_0), .d0(n1423), .sl(net149681), .d1(n1424) );
	inv_16 U2179 ( .x(n866), .a(n865) );
	mux2i_1 U218 ( .x(n3893), .d0(n1680), .sl(n1650), .d1(n1343) );
	inv_2 U2180 ( .x(n868), .a(n1493) );
	nand2i_0 U2181 ( .x(n1493), .a(n1688), .b(n1468) );
	mux2i_1 U2182 ( .x(___cell__36997_net129654), .d0(n2632), .sl(n738), .d1(n1471) );
	buf_16 U2184 ( .x(Imm[20]), .a(N6368) );
	buf_16 U2185 ( .x(Imm[11]), .a(N6350) );
	buf_8 U2186 ( .x(n889), .a(n338) );
	mux2i_8 U2187 ( .x(n339), .d0(n1332), .sl(net149681), .d1(n1333) );
	mux2i_3 U2189 ( .x(reg_dst_of_EX_0), .d0(n561), .sl(reg_dst), .d1(n669) );
	mux2i_1 U219 ( .x(n3897), .d0(n1676), .sl(n1650), .d1(n1338) );
	mux2i_3 U2190 ( .x(reg_dst_of_EX_4), .d0(n558), .sl(reg_dst), .d1(n562) );
	inv_5 U2192 ( .x(n882), .a(n1433) );
	nand2i_2 U2193 ( .x(n1433), .a(CLI), .b(INT) );
	nand2_0 U2194 ( .x(n1717), .a(n642), .b(reg_dst) );
	inv_0 U2196 ( .x(n1543), .a(NPC[11]) );
	aoi222_1 U2197 ( .x(n999), .a(n726), .b(n1719), .c(n1732), .d(EPC_11),
		.e(Cause_Reg_11), .f(n1803) );
	mux2i_1 U2199 ( .x(IR_latched_15), .d0(n568), .sl(net149680), .d1(n1412) );
	nor3_1 U22 ( .x(n1579), .a(n3923), .b(opcode_of_MEM_3), .c(opcode_of_MEM_4) );
	inv_2 U220 ( .x(n1676), .a(N510) );
	inv_0 U2200 ( .x(n1063), .a(n887) );
	oai21_1 U2201 ( .x(N6744), .a(___cell__36997_net125989), .b(n1777), .c(n1023) );
	nand2i_2 U2202 ( .x(___cell__36997_net129657), .a(n1495), .b(n867) );
	nand2i_2 U2203 ( .x(n1146), .a(n1500), .b(n863) );
	nand2i_2 U2204 ( .x(n1187), .a(n1503), .b(n862) );
	nand2i_2 U2205 ( .x(n1199), .a(n1504), .b(n863) );
	nand2i_2 U2206 ( .x(n1251), .a(n1502), .b(n862) );
	aoi21_1 U2208 ( .x(n1180), .a(N5368), .b(n863), .c(n1297) );
	aoi21_1 U2209 ( .x(n1188), .a(N5362), .b(n863), .c(n1300) );
	nand2i_2 U2210 ( .x(n1195), .a(n1506), .b(n862) );
	aoi21_1 U2211 ( .x(n1156), .a(N5351), .b(n863), .c(n1301) );
	nand2i_2 U2213 ( .x(n1234), .a(n1509), .b(n863) );
	aoi21_3 U2214 ( .x(n1256), .a(N5353), .b(n862), .c(n1293) );
	aoi21_3 U2215 ( .x(n1241), .a(N5354), .b(n863), .c(n1275) );
	aoi22_1 U2217 ( .x(n1168), .a(N5359), .b(n895), .c(N6026), .d(___cell__36997_net130214) );
	aoi22_1 U2218 ( .x(n1160), .a(N5367), .b(n895), .c(N6034), .d(___cell__36997_net130214) );
	aoi22_1 U2219 ( .x(n1224), .a(N5363), .b(n895), .c(N6030), .d(___cell__36997_net130214) );
	mux2i_1 U222 ( .x(n1090), .d0(n1587), .sl(___cell__36997_net126612), .d1(n883) );
	aoi22_1 U2221 ( .x(n1151), .a(N5371), .b(n895), .c(N6038), .d(___cell__36997_net130214) );
	oai21_1 U2222 ( .x(n3801), .a(n1053), .b(n3995), .c(n1054) );
	oai21_1 U2223 ( .x(n3775), .a(n725), .b(n1065), .c(n1110) );
	inv_0 U2224 ( .x(n1545), .a(NPC[9]) );
	aoi222_1 U2225 ( .x(n1033), .a(n746), .b(n1719), .c(n1732), .d(EPC_9),
		.e(Cause_Reg_9), .f(n1803) );
	mux2i_1 U2226 ( .x(IR_latched_5), .d0(n565), .sl(n731), .d1(n1417) );
	oai21_1 U2227 ( .x(N6745), .a(n1024), .b(n678), .c(n1025) );
	inv_0 U2228 ( .x(n1547), .a(NPC[7]) );
	aoi222_1 U2229 ( .x(n1243), .a(n554), .b(n1719), .c(n1732), .d(EPC_7),
		.e(Cause_Reg_7), .f(n1803) );
	mux2i_1 U223 ( .x(n3910), .d0(n1663), .sl(n1650), .d1(n1400) );
	inv_0 U2230 ( .x(n1542), .a(NPC[12]) );
	aoi222_1 U2231 ( .x(n1002), .a(NPC[12]), .b(n1802), .c(n1732), .d(EPC_12),
		.e(Cause_Reg_12), .f(n1803) );
	buf_16 U2232 ( .x(reg_out_A[24]), .a(n3957) );
	exor2_1 U2233 ( .x(n1568), .a(IR_opcode_field[2]), .b(IR_opcode_field[4]) );
	nand2i_2 U2234 ( .x(n3812), .a(n1118), .b(n763) );
	buf_16 U2235 ( .x(Imm[28]), .a(N6384) );
	oai21_1 U2236 ( .x(N6743), .a(n698), .b(n995), .c(n1022) );
	nand2i_2 U2237 ( .x(n3809), .a(n1120), .b(n1100) );
	oai21_1 U2238 ( .x(n3802), .a(n1055), .b(n854), .c(n1056) );
	inv_0 U2239 ( .x(n1548), .a(NPC[5]) );
	inv_2 U224 ( .x(n1663), .a(N523) );
	aoi222_1 U2240 ( .x(n1126), .a(n717), .b(n1802), .c(n1732), .d(EPC_5),
		.e(Cause_Reg_5), .f(n1803) );
	inv_7 U2242 ( .x(net148915), .a(___cell__36997_net130217) );
	nand2_0 U2243 ( .x(n1112), .a(n1718), .b(IR_opcode_field[3]) );
	inv_0 U2244 ( .x(n1322), .a(IR_opcode_field[3]) );
	nor2_0 U2245 ( .x(n1700), .a(IR_opcode_field[3]), .b(IR_opcode_field[4]) );
	nand4i_1 U2247 ( .x(n1773), .a(n1734), .b(n1572), .c(n1735), .d(n1444) );
	oai21_1 U2248 ( .x(n3787), .a(n1071), .b(n1775), .c(n1072) );
	exor2_1 U2249 ( .x(n1687), .a(n1686), .b(n1071) );
	buf_16 U2250 ( .x(Imm[17]), .a(N6362) );
	buf_16 U2251 ( .x(Imm[15]), .a(N6358) );
	aoi221_1 U2252 ( .x(n1232), .a(N5440), .b(___cell__36997_net130212), .c(branch_address[21]),
		.d(net148865), .e(n1290) );
	aoi221_1 U2253 ( .x(n1193), .a(N5442), .b(___cell__36997_net130212), .c(branch_address[23]),
		.d(net148865), .e(n1286) );
	aoi22_1 U2254 ( .x(n1162), .a(branch_address[16]), .b(net148865), .c(N5435),
		.d(___cell__36997_net130212) );
	aoi22_1 U2255 ( .x(n1158), .a(branch_address[0]), .b(net148865), .c(N5419),
		.d(___cell__36997_net130212) );
	aoi22_1 U2256 ( .x(n1166), .a(branch_address[14]), .b(net148865), .c(N5433),
		.d(___cell__36997_net130212) );
	aoi22_1 U2257 ( .x(n1170), .a(branch_address[8]), .b(net148865), .c(N5427),
		.d(___cell__36997_net130212) );
	aoi22_1 U2258 ( .x(n1230), .a(branch_address[10]), .b(net148865), .c(N5429),
		.d(___cell__36997_net130212) );
	aoi22_1 U2259 ( .x(n1206), .a(branch_address[9]), .b(net148865), .c(N5428),
		.d(___cell__36997_net130709) );
	mux2i_1 U226 ( .x(n3900), .d0(n1673), .sl(n1650), .d1(n1374) );
	aoi22_1 U2260 ( .x(n1226), .a(branch_address[12]), .b(net148865), .c(N5431),
		.d(___cell__36997_net130212) );
	aoi22_1 U2261 ( .x(n1202), .a(branch_address[4]), .b(net148865), .c(N5423),
		.d(___cell__36997_net130212) );
	aoi22_1 U2262 ( .x(n1221), .a(branch_address[18]), .b(net148865), .c(N5437),
		.d(___cell__36997_net130212) );
	aoi22_1 U2263 ( .x(n1185), .a(branch_address[25]), .b(net148865), .c(n1336),
		.d(n797) );
	buf_16 U2265 ( .x(reg_out_A[7]), .a(n3971) );
	buf_16 U2266 ( .x(reg_out_A[3]), .a(n3974) );
	buf_16 U2267 ( .x(reg_out_A[16]), .a(n3965) );
	buf_16 U2268 ( .x(reg_out_A[8]), .a(n3970) );
	buf_16 U2269 ( .x(Imm[2]), .a(N6332) );
	inv_2 U227 ( .x(n1673), .a(N513) );
	buf_16 U2270 ( .x(Imm[4]), .a(N6336) );
	buf_16 U2271 ( .x(reg_out_A[17]), .a(n3964) );
	nand2_2 U2272 ( .x(n2641), .a(___cell__36997_net126604), .b(n1034) );
	nand2i_4 U2273 ( .x(n3807), .a(n1099), .b(n763) );
	nand2i_4 U2274 ( .x(n3813), .a(n1103), .b(n764) );
	nand2i_4 U2275 ( .x(n3822), .a(n1105), .b(n764) );
	nand2i_4 U2276 ( .x(n3820), .a(n1115), .b(n764) );
	nand2i_4 U2277 ( .x(n3821), .a(n1116), .b(n764) );
	nand2i_4 U2278 ( .x(n3818), .a(n1117), .b(n764) );
	nand2i_4 U2279 ( .x(n3816), .a(n1119), .b(n763) );
	inv_2 U228 ( .x(n1249), .a(n733) );
	nand2i_4 U2280 ( .x(n3819), .a(n1121), .b(n763) );
	nand2i_4 U2281 ( .x(n3808), .a(n1123), .b(n763) );
	nand2i_4 U2282 ( .x(n3817), .a(n1124), .b(n763) );
	nand2i_4 U2283 ( .x(n3814), .a(n1125), .b(n1100) );
	nand4_1 U2284 ( .x(n3851), .a(n1144), .b(n1147), .c(n1146), .d(n1145) );
	nand4_1 U2285 ( .x(n3844), .a(n1151), .b(n1149), .c(n1150), .d(n1148) );
	nand4_1 U2286 ( .x(n3825), .a(n1152), .b(n1153), .c(n1154), .d(n1155) );
	nand4_1 U2287 ( .x(n3824), .a(n1156), .b(n1157), .c(n1158), .d(n1159) );
	nand4_1 U2288 ( .x(n3840), .a(n1160), .b(n1161), .c(n1162), .d(n1163) );
	nand4_1 U2289 ( .x(n3838), .a(n1164), .b(n1165), .c(n1166), .d(n1167) );
	inv_2 U229 ( .x(n1501), .a(N6044) );
	nand4_1 U2290 ( .x(n3832), .a(n1168), .b(n1169), .c(n1170), .d(n1171) );
	nand4_1 U2291 ( .x(n3829), .a(n1172), .b(n1173), .c(n1174), .d(n1175) );
	nand4_1 U2293 ( .x(n3841), .a(n1180), .b(n1181), .c(n1182), .d(n1183) );
	nand4_1 U2294 ( .x(n3835), .a(n1188), .b(n1189), .c(n1190), .d(n1191) );
	nand4_1 U2296 ( .x(n3828), .a(n1200), .b(n1201), .c(n1202), .d(n1203) );
	nand4_1 U2297 ( .x(n3833), .a(n1204), .b(n1206), .c(n1207), .d(n1205) );
	nand4_1 U2298 ( .x(n3843), .a(n1208), .b(n1210), .c(n1209), .d(n1211) );
	nand4_1 U2299 ( .x(n3837), .a(n1212), .b(n1213), .c(n1214), .d(n1215) );
	oa21_2 U23 ( .x(n3923), .a(opcode_of_MEM_2), .b(n3924), .c(opcode_of_MEM_1) );
	inv_2 U230 ( .x(n1502), .a(N5377) );
	nand4_1 U2300 ( .x(n3839), .a(n1218), .b(n1217), .c(n1216), .d(n1219) );
	nand4_1 U2301 ( .x(n3836), .a(n1224), .b(n1225), .c(n1226), .d(n1227) );
	nand4_1 U2302 ( .x(n3834), .a(n1228), .b(n1229), .c(n1230), .d(n1231) );
	nand4_1 U2304 ( .x(n3831), .a(n1246), .b(n1244), .c(n1245), .d(n1247) );
	nand4_1 U2305 ( .x(n3850), .a(n1248), .b(n1249), .c(n1250), .d(n1251) );
	nor2_5 U2306 ( .x(n1184), .a(___cell__36997_net129247), .b(n1281) );
	nor2_5 U2307 ( .x(n1254), .a(___cell__36997_net129247), .b(n1292) );
	nor2_5 U2308 ( .x(n1220), .a(n1272), .b(n1296) );
	nor2_5 U2309 ( .x(n1119), .a(n705), .b(n816) );
	mux2i_1 U231 ( .x(n3895), .d0(n1678), .sl(n1650), .d1(n1346) );
	nor2_5 U2310 ( .x(n1125), .a(n705), .b(n827) );
	nor2_5 U2311 ( .x(n1103), .a(n1776), .b(n789) );
	nor2_5 U2312 ( .x(n1118), .a(n705), .b(n649) );
	nor2_5 U2313 ( .x(n1123), .a(n705), .b(n803) );
	nor2_5 U2314 ( .x(n1099), .a(n1776), .b(n648) );
	mux2i_3 U2315 ( .x(n1258), .d0(n567), .sl(net149680), .d1(n1331) );
	mux2i_3 U2316 ( .x(n1344), .d0(n1345), .sl(___cell__36997_net129354), .d1(n1346) );
	mux2i_3 U2317 ( .x(n1350), .d0(n1351), .sl(___cell__36997_net129354), .d1(n1304) );
	mux2i_3 U2318 ( .x(n1352), .d0(n1353), .sl(___cell__36997_net129354), .d1(n1354) );
	mux2i_3 U2319 ( .x(___cell__36997_net129378), .d0(n1358), .sl(___cell__36997_net129354),
		.d1(n1359) );
	inv_2 U232 ( .x(n1678), .a(N508) );
	mux2i_3 U2320 ( .x(___cell__36997_net129381), .d0(n1360), .sl(___cell__36997_net129354),
		.d1(n1361) );
	mux2i_3 U2321 ( .x(n1364), .d0(n1365), .sl(___cell__36997_net129354), .d1(n1366) );
	mux2i_3 U2322 ( .x(n1369), .d0(n1370), .sl(___cell__36997_net129354), .d1(n1371) );
	mux2i_3 U2323 ( .x(n1372), .d0(n1373), .sl(___cell__36997_net129354), .d1(n1374) );
	mux2i_3 U2324 ( .x(n1388), .d0(n1389), .sl(___cell__36997_net129354), .d1(n1390) );
	mux2i_3 U2325 ( .x(n1393), .d0(n1394), .sl(___cell__36997_net129354), .d1(n1395) );
	mux2i_3 U2326 ( .x(n1398), .d0(n1399), .sl(___cell__36997_net129354), .d1(n1400) );
	mux2i_3 U2327 ( .x(n1401), .d0(n1402), .sl(___cell__36997_net129354), .d1(n1403) );
	mux2i_3 U2328 ( .x(n1404), .d0(n1405), .sl(___cell__36997_net129354), .d1(n1406) );
	mux2i_3 U2329 ( .x(n1407), .d0(n1408), .sl(___cell__36997_net129354), .d1(n1409) );
	mux2i_1 U233 ( .x(n3915), .d0(n1658), .sl(n1650), .d1(n1385) );
	mux2i_3 U2330 ( .x(IR_latched_14), .d0(n569), .sl(net149681), .d1(n1413) );
	mux2i_3 U2331 ( .x(IR_latched_13), .d0(n570), .sl(net149680), .d1(n1414) );
	mux2i_3 U2332 ( .x(IR_latched_11), .d0(n571), .sl(net149680), .d1(n1416) );
	mux2i_3 U2333 ( .x(n1051), .d0(current_IR_9), .sl(net149680), .d1(IR_latched_input[9]) );
	mux2i_3 U2334 ( .x(n1049), .d0(current_IR_8), .sl(n728), .d1(IR_latched_input[8]) );
	oai21_4 U2335 ( .x(n1451), .a(n1450), .b(n556), .c(n1452) );
	oai21_4 U2336 ( .x(n1476), .a(n1477), .b(n1478), .c(n1475) );
	nand2i_4 U2337 ( .x(n1108), .a(n1486), .b(n1430) );
	inv_6 U2338 ( .x(n1419), .a(IR_latched_input[4]) );
	inv_6 U2339 ( .x(n1273), .a(N5381) );
	inv_2 U234 ( .x(n1658), .a(N528) );
	inv_6 U2340 ( .x(n1505), .a(N6042) );
	inv_6 U2341 ( .x(n1296), .a(N5369) );
	exor2_3 U2342 ( .x(n1563), .a(reg_dst_of_MEM_0), .b(n879) );
	exor2_3 U2343 ( .x(n1457), .a(reg_dst_of_MEM_4), .b(n1132) );
	exor2_3 U2344 ( .x(n1569), .a(WB_index_2), .b(n1426) );
	exor2_3 U2345 ( .x(n1572), .a(WB_index_4), .b(n1132) );
	inv_6 U2346 ( .x(n1345), .a(N441) );
	inv_6 U2347 ( .x(n1348), .a(N451) );
	inv_6 U2348 ( .x(n1351), .a(N453) );
	inv_6 U2349 ( .x(n1353), .a(N457) );
	mux2i_1 U235 ( .x(n3751), .d0(n657), .sl(___cell__36997_net130681), .d1(n1329) );
	inv_6 U2350 ( .x(n1358), .a(N454) );
	inv_6 U2351 ( .x(n1360), .a(N442) );
	inv_6 U2354 ( .x(n1370), .a(N467) );
	inv_6 U2355 ( .x(n1373), .a(N446) );
	inv_6 U2356 ( .x(n1378), .a(N447) );
	inv_6 U2357 ( .x(n1384), .a(N461) );
	inv_6 U2358 ( .x(n1389), .a(N466) );
	inv_6 U2359 ( .x(n1394), .a(N460) );
	aoi222_1 U236 ( .x(n1023), .a(NPC[26]), .b(n1802), .c(n1732), .d(EPC_26),
		.e(Cause_Reg_26), .f(n1803) );
	inv_6 U2360 ( .x(n1405), .a(N455) );
	inv_6 U2361 ( .x(n1408), .a(N444) );
	mux2i_3 U2362 ( .x(n3761), .d0(n656), .sl(___cell__36997_net126612), .d1(n3992) );
	mux2i_3 U2363 ( .x(n3421), .d0(n2630), .sl(n1857), .d1(n1800) );
	mux2i_3 U2364 ( .x(n3444), .d0(n2629), .sl(n1857), .d1(n1799) );
	mux2i_3 U2365 ( .x(n3453), .d0(n2606), .sl(n1856), .d1(n1603) );
	mux2i_3 U2366 ( .x(n3476), .d0(n2605), .sl(n1856), .d1(n1799) );
	mux2i_3 U2367 ( .x(n3485), .d0(n2582), .sl(n1855), .d1(n1800) );
	mux2i_3 U2368 ( .x(n3508), .d0(n2581), .sl(n1855), .d1(n1799) );
	mux2i_3 U2369 ( .x(n3517), .d0(n2558), .sl(n1854), .d1(n1603) );
	aoi22_2 U237 ( .x(n1148), .a(branch_address[20]), .b(n766), .c(N5439),
		.d(___cell__36997_net130212) );
	mux2i_3 U2370 ( .x(n3540), .d0(n2557), .sl(n1854), .d1(n1799) );
	mux2i_3 U2371 ( .x(n3549), .d0(n2534), .sl(n1853), .d1(n1800) );
	mux2i_3 U2372 ( .x(n3572), .d0(n2533), .sl(n1853), .d1(n1799) );
	mux2i_3 U2373 ( .x(n3581), .d0(n2510), .sl(n1852), .d1(n1603) );
	mux2i_3 U2374 ( .x(n3604), .d0(n2509), .sl(n1852), .d1(n1799) );
	mux2i_3 U2375 ( .x(n3613), .d0(n2486), .sl(n1851), .d1(n1800) );
	mux2i_3 U2376 ( .x(n3636), .d0(n2485), .sl(n1851), .d1(n1799) );
	mux2i_3 U2377 ( .x(n2717), .d0(n2462), .sl(n1850), .d1(n1603) );
	mux2i_3 U2378 ( .x(n2740), .d0(n2461), .sl(n1850), .d1(n1799) );
	mux2i_3 U2379 ( .x(n2749), .d0(n2438), .sl(n1849), .d1(n1800) );
	mux2i_1 U238 ( .x(n3904), .d0(n1669), .sl(n1650), .d1(n1340) );
	mux2i_3 U2380 ( .x(n2772), .d0(n2437), .sl(n1849), .d1(n1799) );
	mux2i_3 U2381 ( .x(n3645), .d0(n2414), .sl(n1848), .d1(n1603) );
	mux2i_3 U2382 ( .x(n3668), .d0(n2413), .sl(n1848), .d1(n1799) );
	mux2i_3 U2383 ( .x(n2781), .d0(n2390), .sl(n1847), .d1(n1800) );
	mux2i_3 U2384 ( .x(n2804), .d0(n2389), .sl(n1847), .d1(n1799) );
	mux2i_3 U2385 ( .x(n2813), .d0(n2366), .sl(n1846), .d1(n1603) );
	mux2i_3 U2386 ( .x(n2836), .d0(n2365), .sl(n1846), .d1(n1799) );
	mux2i_3 U2387 ( .x(n2845), .d0(n2342), .sl(n1845), .d1(n1800) );
	mux2i_3 U2388 ( .x(n2868), .d0(n2341), .sl(n1845), .d1(n1799) );
	mux2i_3 U2389 ( .x(n2877), .d0(n2318), .sl(n1844), .d1(n1603) );
	inv_2 U239 ( .x(n1669), .a(N517) );
	mux2i_3 U2390 ( .x(n2900), .d0(n2317), .sl(n1844), .d1(n1799) );
	mux2i_3 U2391 ( .x(n2909), .d0(n2294), .sl(n1843), .d1(n1800) );
	mux2i_3 U2392 ( .x(n2932), .d0(n2293), .sl(n1843), .d1(n1799) );
	mux2i_3 U2393 ( .x(n2941), .d0(n2270), .sl(n1842), .d1(n1603) );
	mux2i_3 U2394 ( .x(n2964), .d0(n2269), .sl(n1842), .d1(n1799) );
	mux2i_3 U2395 ( .x(n2973), .d0(n2246), .sl(n1841), .d1(n1603) );
	mux2i_3 U2396 ( .x(n2996), .d0(n2245), .sl(n1841), .d1(n1799) );
	mux2i_3 U2397 ( .x(n3005), .d0(n2222), .sl(n1840), .d1(n1800) );
	mux2i_3 U2398 ( .x(n3028), .d0(n2221), .sl(n1840), .d1(n1799) );
	mux2i_3 U2399 ( .x(n3037), .d0(n2198), .sl(n1839), .d1(n1603) );
	nand2_2 U24 ( .x(n3946), .a(n3945), .b(n3924) );
	mux2i_1 U240 ( .x(n3909), .d0(n1664), .sl(n1650), .d1(n1406) );
	mux2i_3 U2400 ( .x(n3060), .d0(n2197), .sl(n1839), .d1(n1799) );
	mux2i_3 U2401 ( .x(n3069), .d0(n2174), .sl(n1838), .d1(n1800) );
	mux2i_3 U2402 ( .x(n3092), .d0(n2173), .sl(n1838), .d1(n1799) );
	mux2i_3 U2403 ( .x(n3677), .d0(n2150), .sl(n1837), .d1(n1800) );
	mux2i_3 U2404 ( .x(n3700), .d0(n2149), .sl(n1837), .d1(n1799) );
	mux2i_3 U2405 ( .x(n3101), .d0(n2126), .sl(n1836), .d1(n1603) );
	mux2i_3 U2406 ( .x(n3124), .d0(n2125), .sl(n1836), .d1(n1799) );
	mux2i_3 U2407 ( .x(n3133), .d0(n2102), .sl(n1835), .d1(n1800) );
	mux2i_3 U2408 ( .x(n3156), .d0(n2101), .sl(n1835), .d1(n1799) );
	mux2i_3 U2409 ( .x(n3165), .d0(n2078), .sl(n1834), .d1(n1603) );
	inv_2 U241 ( .x(n1664), .a(N522) );
	mux2i_3 U2410 ( .x(n3188), .d0(n2077), .sl(n1834), .d1(n1799) );
	mux2i_3 U2411 ( .x(n3197), .d0(n2054), .sl(n1833), .d1(n1800) );
	mux2i_3 U2412 ( .x(n3220), .d0(n2053), .sl(n1833), .d1(n1799) );
	mux2i_3 U2413 ( .x(n3229), .d0(n2030), .sl(n1832), .d1(n1603) );
	mux2i_3 U2414 ( .x(n3252), .d0(n2029), .sl(n1832), .d1(n1799) );
	mux2i_3 U2415 ( .x(n3261), .d0(n2006), .sl(n1831), .d1(n1800) );
	mux2i_3 U2416 ( .x(n3284), .d0(n2005), .sl(n1831), .d1(n1799) );
	mux2i_3 U2417 ( .x(n3293), .d0(n1982), .sl(n1830), .d1(n1603) );
	mux2i_3 U2418 ( .x(n3316), .d0(n1981), .sl(n1830), .d1(n1799) );
	mux2i_3 U2419 ( .x(n3325), .d0(n1958), .sl(n1829), .d1(n1603) );
	mux2i_3 U2420 ( .x(n3348), .d0(n1957), .sl(n1829), .d1(n1799) );
	mux2i_3 U2421 ( .x(n3357), .d0(n1934), .sl(n1828), .d1(n1800) );
	mux2i_3 U2422 ( .x(n3380), .d0(n1933), .sl(n1828), .d1(n1799) );
	mux2i_3 U2423 ( .x(n3389), .d0(n1910), .sl(n1827), .d1(n1800) );
	mux2i_3 U2424 ( .x(n3412), .d0(n1909), .sl(n1827), .d1(n1799) );
	mux2i_3 U2425 ( .x(n3710), .d0(n1887), .sl(n1826), .d1(n1801) );
	mux2i_3 U2426 ( .x(n3709), .d0(n1886), .sl(n1826), .d1(n1603) );
	mux2i_3 U2427 ( .x(n3732), .d0(n1885), .sl(n1826), .d1(n1799) );
	mux2i_3 U2428 ( .x(n3731), .d0(n1884), .sl(n1826), .d1(n1798) );
	mux2i_3 U2429 ( .x(n3730), .d0(n1883), .sl(n1826), .d1(n1797) );
	nand2i_2 U243 ( .x(n1046), .a(n643), .b(n1718) );
	mux2i_3 U2430 ( .x(n3729), .d0(n1882), .sl(n1826), .d1(n1796) );
	mux2i_3 U2431 ( .x(n3728), .d0(n1881), .sl(n1826), .d1(n1795) );
	mux2i_3 U2432 ( .x(n3727), .d0(n1880), .sl(n1826), .d1(n1794) );
	mux2i_3 U2433 ( .x(n3726), .d0(n1879), .sl(n1826), .d1(n1793) );
	mux2i_3 U2434 ( .x(n3725), .d0(n1878), .sl(n1826), .d1(n1792) );
	mux2i_3 U2435 ( .x(n3724), .d0(n1877), .sl(n1826), .d1(n1791) );
	mux2i_3 U2436 ( .x(n3723), .d0(n1876), .sl(n1826), .d1(n1790) );
	mux2i_3 U2437 ( .x(n3722), .d0(n1875), .sl(n1826), .d1(n1789) );
	mux2i_3 U2438 ( .x(n3721), .d0(n1874), .sl(n1826), .d1(n1788) );
	mux2i_3 U2439 ( .x(n3720), .d0(n1873), .sl(n1826), .d1(n1787) );
	mux2i_3 U2440 ( .x(n3719), .d0(n1872), .sl(n1826), .d1(n1786) );
	mux2i_3 U2441 ( .x(n3718), .d0(n1871), .sl(n1826), .d1(n1785) );
	mux2i_3 U2442 ( .x(n3717), .d0(n1870), .sl(n1826), .d1(n1784) );
	mux2i_3 U2443 ( .x(n3716), .d0(n1869), .sl(n1826), .d1(n1783) );
	mux2i_3 U2444 ( .x(n3715), .d0(n1868), .sl(n1826), .d1(n1782) );
	mux2i_3 U2445 ( .x(n3714), .d0(n1867), .sl(n1826), .d1(n1781) );
	mux2i_3 U2446 ( .x(n3713), .d0(n1866), .sl(n1826), .d1(n1780) );
	mux2i_3 U2447 ( .x(n3712), .d0(n1865), .sl(n1826), .d1(n1779) );
	mux2i_3 U2448 ( .x(n3711), .d0(n1864), .sl(n1826), .d1(n1778) );
	mux2i_3 U2449 ( .x(n2651), .d0(n618), .sl(___cell__36997_net130567), .d1(n873) );
	nand2i_2 U245 ( .x(n1048), .a(n734), .b(n642) );
	mux2i_3 U2450 ( .x(n2650), .d0(n619), .sl(___cell__36997_net130125), .d1(n872) );
	mux2i_3 U2451 ( .x(n2649), .d0(n620), .sl(___cell__36997_net130567), .d1(n734) );
	mux2i_3 U2452 ( .x(n2648), .d0(n621), .sl(___cell__36997_net130125), .d1(n643) );
	mux2i_3 U2453 ( .x(n2672), .d0(n597), .sl(___cell__36997_net130125), .d1(n701) );
	mux2i_3 U2454 ( .x(n2645), .d0(n624), .sl(___cell__36997_net130567), .d1(n886) );
	mux2i_3 U2455 ( .x(n2671), .d0(n598), .sl(___cell__36997_net130125), .d1(n762) );
	mux2i_3 U2456 ( .x(n2670), .d0(n599), .sl(___cell__36997_net130567), .d1(n696) );
	mux2i_3 U2457 ( .x(n2669), .d0(n600), .sl(___cell__36997_net130125), .d1(n765) );
	mux2i_3 U2458 ( .x(n2668), .d0(n601), .sl(___cell__36997_net130567), .d1(n735) );
	mux2i_3 U2459 ( .x(n2667), .d0(n602), .sl(___cell__36997_net130125), .d1(n816) );
	mux2i_3 U2460 ( .x(n2665), .d0(n604), .sl(___cell__36997_net130125), .d1(n827) );
	mux2i_3 U2461 ( .x(n2664), .d0(n605), .sl(___cell__36997_net130567), .d1(n789) );
	mux2i_3 U2462 ( .x(n2663), .d0(n606), .sl(___cell__36997_net130125), .d1(n649) );
	mux2i_3 U2463 ( .x(n2662), .d0(n607), .sl(___cell__36997_net130567), .d1(n732) );
	mux2i_3 U2464 ( .x(n2644), .d0(n625), .sl(___cell__36997_net130125), .d1(n870) );
	mux2i_3 U2465 ( .x(n2661), .d0(n608), .sl(___cell__36997_net130567), .d1(n775) );
	mux2i_3 U2466 ( .x(n2660), .d0(n609), .sl(___cell__36997_net130125), .d1(n778) );
	mux2i_3 U2467 ( .x(n2659), .d0(n610), .sl(___cell__36997_net130567), .d1(n803) );
	mux2i_3 U2468 ( .x(n2658), .d0(n611), .sl(___cell__36997_net130125), .d1(n648) );
	mux2i_3 U2469 ( .x(n2657), .d0(n612), .sl(___cell__36997_net130567), .d1(n829) );
	nand2i_4 U247 ( .x(n1058), .a(n779), .b(n642) );
	mux2i_3 U2470 ( .x(n2656), .d0(n613), .sl(___cell__36997_net130125), .d1(n647) );
	mux2i_3 U2471 ( .x(n2654), .d0(n615), .sl(___cell__36997_net130125), .d1(n779) );
	mux2i_3 U2472 ( .x(n2653), .d0(n616), .sl(___cell__36997_net130567), .d1(n786) );
	mux2i_3 U2473 ( .x(n2643), .d0(n626), .sl(___cell__36997_net130567), .d1(n720) );
	nand4_1 U2474 ( .x(n1486), .a(n739), .b(n1081), .c(n1067), .d(n767) );
	and4i_5 U2475 ( .x(n1447), .a(n1558), .b(n1697), .c(n1696), .d(n1695) );
	and3i_4 U2477 ( .x(___cell__36997_net130187), .a(n1685), .b(reg_write_WB),
		.c(n1569) );
	nor2_5 U2478 ( .x(n1705), .a(___cell__36997_net130191), .b(n1704) );
	nor2_5 U2479 ( .x(n1708), .a(n1706), .b(n1707) );
	mux2i_1 U248 ( .x(n3903), .d0(n1670), .sl(n1650), .d1(n1383) );
	nor2_5 U2480 ( .x(n1711), .a(n1709), .b(n1710) );
	inv_6 U2481 ( .x(n1654), .a(N531) );
	inv_5 U2482 ( .x(n1857), .a(n1741) );
	inv_5 U2483 ( .x(n1856), .a(n1742) );
	inv_5 U2484 ( .x(n1855), .a(n1743) );
	inv_5 U2485 ( .x(n1854), .a(n1744) );
	inv_5 U2486 ( .x(n1853), .a(n1745) );
	inv_5 U2487 ( .x(n1852), .a(n1746) );
	inv_5 U2488 ( .x(n1851), .a(n1747) );
	inv_5 U2489 ( .x(n1850), .a(n1748) );
	inv_2 U249 ( .x(n1670), .a(N516) );
	inv_5 U2490 ( .x(n1849), .a(n1749) );
	inv_5 U2491 ( .x(n1848), .a(n1750) );
	inv_5 U2492 ( .x(n1847), .a(n1751) );
	inv_5 U2493 ( .x(n1846), .a(n1752) );
	inv_5 U2494 ( .x(n1845), .a(n1753) );
	inv_5 U2495 ( .x(n1844), .a(n1754) );
	inv_5 U2496 ( .x(n1843), .a(n1755) );
	inv_5 U2497 ( .x(n1842), .a(n1756) );
	inv_5 U2498 ( .x(n1841), .a(n1757) );
	inv_5 U2499 ( .x(n1840), .a(n1758) );
	nand2_2 U25 ( .x(n3947), .a(n556), .b(n3932) );
	mux2i_1 U250 ( .x(n3908), .d0(n1665), .sl(n1650), .d1(n1359) );
	inv_5 U2500 ( .x(n1839), .a(n1759) );
	inv_5 U2501 ( .x(n1838), .a(n1760) );
	inv_5 U2502 ( .x(n1837), .a(n1761) );
	inv_5 U2503 ( .x(n1836), .a(n1762) );
	inv_5 U2504 ( .x(n1835), .a(n1763) );
	inv_5 U2505 ( .x(n1834), .a(n1764) );
	inv_5 U2506 ( .x(n1833), .a(n1765) );
	inv_5 U2507 ( .x(n1832), .a(n1766) );
	inv_5 U2508 ( .x(n1831), .a(n1767) );
	inv_5 U2509 ( .x(n1830), .a(n1768) );
	inv_2 U251 ( .x(n1665), .a(N521) );
	inv_5 U2510 ( .x(n1829), .a(n1769) );
	inv_5 U2511 ( .x(n1828), .a(n1770) );
	inv_5 U2512 ( .x(n1827), .a(n1771) );
	inv_5 U2513 ( .x(n1826), .a(n1772) );
	buf_16 U2514 ( .x(n331), .a(n761) );
	buf_16 U2515 ( .x(n336), .a(n1258) );
	buf_16 U2516 ( .x(Imm[0]), .a(N6328) );
	buf_16 U2517 ( .x(Imm[5]), .a(N6338) );
	buf_16 U2518 ( .x(Imm[29]), .a(N6386) );
	buf_16 U2519 ( .x(Imm[30]), .a(N6388) );
	mux2i_1 U252 ( .x(n3917), .d0(n1655), .sl(n1650), .d1(n1368) );
	buf_16 U2520 ( .x(reg_out_B[4]), .a(n3980) );
	buf_16 U2521 ( .x(reg_out_B[1]), .a(n3983) );
	buf_16 U2522 ( .x(reg_out_A[4]), .a(n3973) );
	buf_16 U2523 ( .x(reg_out_A[19]), .a(n3962) );
	buf_16 U2524 ( .x(reg_out_A[18]), .a(n3963) );
	buf_16 U2525 ( .x(reg_out_B[3]), .a(n3981) );
	buf_16 U2526 ( .x(reg_out_A[21]), .a(n3960) );
	buf_16 U2527 ( .x(reg_out_A[30]), .a(n3951) );
	nand2i_5 U2528 ( .x(___cell__36997_net126604), .a(___cell__36997_net127190),
		.b(n1484) );
	nand2i_6 U2529 ( .x(n1776), .a(___cell__36997_net130681), .b(n1461) );
	inv_2 U253 ( .x(n1655), .a(N530) );
	nand2i_5 U2531 ( .x(n1145), .a(n1499), .b(___cell__36997_net130212) );
	aoai211_5 U2532 ( .x(n1134), .a(n1570), .b(n1494), .c(n1712), .d(___cell__36997_net126612) );
	nand2i_8 U2533 ( .x(___cell__36997_net127190), .a(n1259), .b(n1461) );
	inv_16 U2534 ( .x(___cell__36997_net126612), .a(___cell__36997_net127190) );
	inv_16 U2535 ( .x(n1132), .a(n336) );
	nand2i_6 U2536 ( .x(___cell__36997_net129626), .a(n1491), .b(n1437) );
	inv_14 U2537 ( .x(n1484), .a(n1471) );
	nand2i_6 U2538 ( .x(n1263), .a(n1470), .b(n860) );
	nand4i_5 U2539 ( .x(n1480), .a(n1264), .b(n1481), .c(n1482), .d(n1483) );
	nand2i_2 U254 ( .x(n1062), .a(n647), .b(n642) );
	inv_14 U2540 ( .x(n1802), .a(n1307) );
	nor2i_8 U2541 ( .x(n1554), .a(n1461), .b(n642) );
	inv_16 U2542 ( .x(n1732), .a(n1518) );
	nand2_8 U2543 ( .x(n1647), .a(n1514), .b(n1648) );
	nand2_8 U2544 ( .x(n1645), .a(n1514), .b(n1646) );
	nand2_8 U2545 ( .x(n1643), .a(n1514), .b(n1644) );
	nand2_8 U2546 ( .x(n1641), .a(n1514), .b(n1642) );
	nand2_8 U2547 ( .x(n1639), .a(n1514), .b(n1640) );
	nand2_8 U2548 ( .x(n1637), .a(n1514), .b(n1638) );
	nand2_8 U2549 ( .x(n1635), .a(n1605), .b(n1636) );
	ao21_1 U255 ( .x(n1473), .a(n1714), .b(___cell__36997_net127190), .c(n1093) );
	nand2_8 U2550 ( .x(n1633), .a(n1605), .b(n1634) );
	nand2_8 U2551 ( .x(n1631), .a(n1605), .b(n1632) );
	nand2_8 U2552 ( .x(n1629), .a(n1605), .b(n1630) );
	nand2_8 U2553 ( .x(n1627), .a(n1605), .b(n1628) );
	nand2_8 U2554 ( .x(n1625), .a(n1605), .b(n1626) );
	nand2_8 U2555 ( .x(n1623), .a(n1605), .b(n1624) );
	nand2_8 U2556 ( .x(n1621), .a(n1605), .b(n1622) );
	nand2_8 U2557 ( .x(n1619), .a(n1605), .b(n1620) );
	nand2_8 U2558 ( .x(n1617), .a(n1605), .b(n1618) );
	nand2_8 U2559 ( .x(n1615), .a(n1605), .b(n1616) );
	inv_5 U256 ( .x(n1494), .a(n1465) );
	nand2_8 U2560 ( .x(n1613), .a(n1605), .b(n1614) );
	nand2_8 U2561 ( .x(n1611), .a(n1605), .b(n1612) );
	nand2_8 U2562 ( .x(n1609), .a(n1605), .b(n1610) );
	nand2_8 U2563 ( .x(n1607), .a(n1605), .b(n1608) );
	nand2_8 U2564 ( .x(n1601), .a(n1514), .b(n1602) );
	inv_16 U2565 ( .x(___cell__36997_net130217), .a(net148858) );
	inv_10 U2566 ( .x(n1492), .a(n1263) );
	nand3_4 U2567 ( .x(n1260), .a(n1460), .b(n564), .c(net152025) );
	nand2_8 U2568 ( .x(n1471), .a(n650), .b(n1436) );
	nand2i_8 U2569 ( .x(n1514), .a(n1723), .b(n1740) );
	mux2i_1 U257 ( .x(n3739), .d0(n1594), .sl(___cell__36997_net130681), .d1(n1595) );
	inv_16 U2570 ( .x(n1605), .a(n1513) );
	nand3i_5 U2571 ( .x(___cell__36997_net129625), .a(n1721), .b(n1465), .c(n834) );
	nand2i_6 U2572 ( .x(n1465), .a(n836), .b(n682) );
	nand2i_8 U2573 ( .x(n1511), .a(N13832), .b(n1512) );
	nand2i_8 U2574 ( .x(n1513), .a(n1302), .b(n1514) );
	nand4_5 U2575 ( .x(n1303), .a(opcode_of_WB_5), .b(n3889), .c(n3887), .d(n3890) );
	exnor2_5 U2577 ( .x(n1558), .a(n1559), .b(n331) );
	exor2_5 U2578 ( .x(n1683), .a(n635), .b(___cell__36997_net129477) );
	mux2i_1 U258 ( .x(n3899), .d0(n1674), .sl(n1650), .d1(n1403) );
	inv_2 U259 ( .x(n1674), .a(N512) );
	exnor2_1 U26 ( .x(n667), .a(reg_dst_of_MEM_1), .b(n1071) );
	mux2i_1 U260 ( .x(n3898), .d0(n1675), .sl(n1650), .d1(n1409) );
	inv_2 U261 ( .x(n1675), .a(N511) );
	inv_2 U2611 ( .x(n1858), .a(reset) );
	inv_2 U2612 ( .x(n848), .a(n1088) );
	inv_7 U2613 ( .x(n749), .a(n3997) );
	inv_7 U2614 ( .x(n1197), .a(n4005) );
	mux2i_1 U2615 ( .x(n815), .d0(n1318), .sl(net149681), .d1(n1319) );
	inv_10 U2616 ( .x(n1081), .a(n712) );
	inv_6 U2617 ( .x(n716), .a(n1317) );
	mux2i_3 U2618 ( .x(n887), .d0(n568), .sl(net149680), .d1(n1412) );
	mux2i_3 U2619 ( .x(n831), .d0(n1418), .sl(net149680), .d1(n1419) );
	mux2i_1 U262 ( .x(n3921), .d0(n1651), .sl(n1650), .d1(n1371) );
	mux2i_6 U2620 ( .x(IR_latched_2), .d0(n1422), .sl(net149236), .d1(n1421) );
	nand4_3 U2621 ( .x(n1709), .a(n1018), .b(n1001), .c(n636), .d(n1031) );
	inv_4 U2622 ( .x(n1367), .a(N463) );
	oa22_3 U2623 ( .x(n823), .a(n724), .b(n711), .c(n1688), .d(n1431) );
	nand4_4 U2624 ( .x(n1707), .a(n638), .b(n1252), .c(n673), .d(n672) );
	nand2_8 U2625 ( .x(___cell__36997_net129624), .a(n1713), .b(n1481) );
	nand2i_5 U2626 ( .x(n1481), .a(n1715), .b(n682) );
	mux2i_3 U2627 ( .x(n3984), .d0(n1376), .sl(n798), .d1(n1375) );
	inv_6 U2628 ( .x(n663), .a(n3984) );
	inv_5 U2629 ( .x(n1375), .a(N452) );
	inv_2 U263 ( .x(n1651), .a(N534) );
	buf_14 U2630 ( .x(net148858), .a(___cell__36997_net127155) );
	inv_6 U2631 ( .x(n799), .a(___cell__36997_net127155) );
	nand4_4 U2632 ( .x(___cell__36997_net130191), .a(n641), .b(___cell__36997_net126005),
		.c(___cell__36997_net125989), .d(___cell__36997_net125941) );
	nand2i_2 U2633 ( .x(n794), .a(n641), .b(n797) );
	inv_0 U2634 ( .x(n3985), .a(n1364) );
	inv_5 U2635 ( .x(n994), .a(n1364) );
	inv_5 U2636 ( .x(n1365), .a(N468) );
	inv_1 U2637 ( .x(n3986), .a(n848) );
	inv_10 U2638 ( .x(n1088), .a(n889) );
	buf_16 U2639 ( .x(reg_out_B[22]), .a(n3977) );
	nand2_2 U264 ( .x(n1114), .a(n642), .b(IR_opcode_field[2]) );
	nand4_1 U2640 ( .x(n3830), .a(n1176), .b(n1177), .c(n1178), .d(n1179) );
	aoi21_4 U2641 ( .x(n1176), .a(N5357), .b(n862), .c(n1269) );
	buf_2 U2642 ( .x(n833), .a(n339) );
	nand3_4 U2643 ( .x(n782), .a(n855), .b(n700), .c(n747) );
	nor3i_2 U2644 ( .x(n1699), .a(n1440), .b(n837), .c(n825) );
	inv_5 U2645 ( .x(n1269), .a(n4007) );
	mux2i_8 U2646 ( .x(n884), .d0(n644), .sl(n736), .d1(IR_latched_input[16]) );
	inv_10 U2647 ( .x(n736), .a(net149236) );
	exnor2_3 U2648 ( .x(n3987), .a(n3988), .b(n879) );
	inv_4 U2649 ( .x(n748), .a(n3987) );
	aoi222_1 U265 ( .x(n1025), .a(NPC[27]), .b(n1719), .c(n1732), .d(EPC_27),
		.e(Cause_Reg_27), .f(n1803) );
	inv_4 U2650 ( .x(n3988), .a(reg_dst_of_EX_0) );
	mux2i_8 U2651 ( .x(n879), .d0(IR_latched_input[21]), .sl(net149236), .d1(current_IR_21) );
	nor2_2 U2652 ( .x(n1464), .a(n1688), .b(n1113) );
	inv_7 U2653 ( .x(n1113), .a(n1315) );
	aoi22_2 U2654 ( .x(n1246), .a(N5426), .b(___cell__36997_net130212), .c(N6025),
		.d(___cell__36997_net130713) );
	aoi211_1 U2655 ( .x(n3989), .a(n1083), .b(n853), .c(n1081), .d(n1113) );
	inv_7 U2656 ( .x(n853), .a(n850) );
	inv_10 U2657 ( .x(n3990), .a(n768) );
	inv_6 U2658 ( .x(n334), .a(n768) );
	buf_10 U2659 ( .x(net149680), .a(___cell__36997_net130572) );
	mux2i_1 U266 ( .x(n3912), .d0(n1661), .sl(n1650), .d1(n1392) );
	buf_14 U2660 ( .x(net149681), .a(n731) );
	buf_4 U2661 ( .x(n837), .a(n1313) );
	nand4_3 U2662 ( .x(n3854), .a(n1135), .b(n758), .c(n1136), .d(n1137) );
	inv_7 U2663 ( .x(n1135), .a(n3996) );
	inv_0 U2664 ( .x(n3991), .a(n1111) );
	inv_2 U2665 ( .x(n3992), .a(n3991) );
	mux2i_6 U2666 ( .x(n1111), .d0(IR_latched_input[29]), .sl(net149236), .d1(current_IR_29) );
	and2_4 U2667 ( .x(n4432), .a(n3910), .b(n681) );
	aoi21_3 U2668 ( .x(n1244), .a(N5358), .b(n863), .c(n1598) );
	inv_6 U2669 ( .x(___cell__36997_net126005), .a(___cell__36997_net129384) );
	inv_2 U267 ( .x(n1661), .a(N525) );
	mux2i_5 U2670 ( .x(___cell__36997_net129384), .d0(n1362), .sl(___cell__36997_net129354),
		.d1(n1363) );
	and4i_3 U2671 ( .x(n1453), .a(n1683), .b(n1698), .c(n1562), .d(n1564) );
	exor2_3 U2672 ( .x(n1564), .a(reg_dst_of_MEM_1), .b(n1565) );
	nand2i_4 U2673 ( .x(n1313), .a(n709), .b(n1453) );
	nand4_3 U2674 ( .x(n3846), .a(n749), .b(n1235), .c(n676), .d(n1236) );
	nand4_3 U2675 ( .x(n3848), .a(n1197), .b(n1196), .c(n1198), .d(n1199) );
	ao22_3 U2676 ( .x(n3993), .a(branch_address[19]), .b(n766), .c(N5438),
		.d(___cell__36997_net130709) );
	inv_4 U2677 ( .x(n1210), .a(n3993) );
	inv_16 U2678 ( .x(___cell__36997_net130709), .a(___cell__36997_net129247) );
	aoi22_3 U2679 ( .x(n1208), .a(N5370), .b(n895), .c(N6037), .d(___cell__36997_net130214) );
	inv_12 U268 ( .x(n724), .a(n739) );
	ao211_5 U2680 ( .x(_branch_address_reg_31_net46811), .a(N5450), .b(n783),
		.c(n664), .d(n792) );
	aoi21_2 U2681 ( .x(n1164), .a(N5365), .b(n862), .c(n1299) );
	nor2i_1 U2682 ( .x(n1299), .a(N6032), .b(___cell__36997_net129239) );
	buf_8 U2683 ( .x(reg_out_B[6]), .a(n4457) );
	aoi21_3 U2684 ( .x(n1139), .a(N5380), .b(n862), .c(n1278) );
	oai21_5 U2685 ( .x(n3995), .a(n1484), .b(n1480), .c(n1554) );
	ao221_5 U2686 ( .x(n3996), .a(___cell__36997_net129384), .b(n797), .c(branch_address[30]),
		.d(n766), .e(n1271) );
	nor2_6 U2687 ( .x(n1271), .a(n1272), .b(n1273) );
	nor2_4 U2688 ( .x(n1286), .a(net148915), .b(n1287) );
	nor2_3 U2689 ( .x(n1295), .a(net148915), .b(n585) );
	inv_2 U269 ( .x(n1504), .a(N5375) );
	inv_5 U2690 ( .x(n1270), .a(n835) );
	ao221_5 U2691 ( .x(n3997), .a(N5441), .b(___cell__36997_net130709), .c(branch_address[22]),
		.d(n766), .e(n1288) );
	nor2_4 U2692 ( .x(n1288), .a(net148913), .b(n1289) );
	inv_16 U2693 ( .x(___cell__36997_net130212), .a(___cell__36997_net129247) );
	inv_3 U2694 ( .x(n1277), .a(N5448) );
	nand4i_2 U2695 ( .x(n3849), .a(n1184), .b(n1186), .c(n1185), .d(n1187) );
	nor2_6 U2696 ( .x(n1290), .a(net148916), .b(n1291) );
	nand4i_1 U2697 ( .x(n792), .a(___cell__36997_net129654), .b(___cell__36997_net129657),
		.c(n794), .d(n793) );
	buf_2 U2698 ( .x(n3998), .a(n805) );
	buf_14 U2699 ( .x(Imm[14]), .a(N6356) );
	buf_14 U27 ( .x(reg_out_A[12]), .a(n3966) );
	inv_2 U270 ( .x(n1510), .a(N6033) );
	buf_14 U2700 ( .x(Imm[6]), .a(N6340) );
	oai22_2 U2701 ( .x(n3795), .a(n705), .b(n871), .c(n3995), .d(n1043) );
	aoi21_2 U2702 ( .x(n1186), .a(N6043), .b(___cell__36997_net130713), .c(n1282) );
	oa22_4 U2703 ( .x(n1204), .a(n4004), .b(n1272), .c(n4003), .d(___cell__36997_net129239) );
	mux2i_8 U2704 ( .x(n3999), .d0(n4001), .sl(n4000), .d1(n4002) );
	inv_0 U2705 ( .x(n1045), .a(n3999) );
	inv_10 U2706 ( .x(n4000), .a(n728) );
	inv_2 U2707 ( .x(n4001), .a(IR_latched_input[6]) );
	inv_2 U2708 ( .x(n4002), .a(current_IR_6) );
	buf_14 U2709 ( .x(n728), .a(n731) );
	nand2i_2 U271 ( .x(n1079), .a(n1861), .b(n642) );
	inv_16 U2710 ( .x(n895), .a(n1272) );
	inv_0 U2711 ( .x(n4003), .a(N6027) );
	inv_0 U2712 ( .x(n4004), .a(N5360) );
	nand2_5 U2713 ( .x(___cell__36997_net129239), .a(net148863), .b(n1494) );
	buf_16 U2714 ( .x(Imm[13]), .a(N6354) );
	buf_8 U2715 ( .x(reg_out_B[2]), .a(n3982) );
	mux2i_8 U2716 ( .x(n817), .d0(n1595), .sl(net152024), .d1(n1594) );
	and2_4 U2717 ( .x(n4442), .a(n3905), .b(n680) );
	inv_8 U2718 ( .x(net148865), .a(n738) );
	ao221_5 U2719 ( .x(n4005), .a(N5443), .b(___cell__36997_net130709), .c(branch_address[24]),
		.d(n766), .e(n1284) );
	nor2_3 U272 ( .x(n1124), .a(n1776), .b(n735) );
	buf_8 U2720 ( .x(n766), .a(n1804) );
	aoi22_2 U2721 ( .x(n1142), .a(branch_address[28]), .b(net148865), .c(N6046),
		.d(___cell__36997_net130214) );
	nor2i_5 U2722 ( .x(n1698), .a(n1563), .b(n1684) );
	buf_10 U2723 ( .x(Imm[16]), .a(N6360) );
	buf_14 U2724 ( .x(Imm[18]), .a(N6364) );
	buf_10 U2725 ( .x(IR_opcode_field[1]), .a(n4453) );
	inv_8 U2726 ( .x(n1130), .a(n1369) );
	nand2i_4 U2727 ( .x(n4007), .a(n4008), .b(___cell__36997_net130214) );
	inv_0 U2728 ( .x(n4008), .a(N6024) );
	exnor2_2 U2729 ( .x(n770), .a(reg_dst_of_EX_1), .b(n339) );
	mux2i_1 U273 ( .x(n3906), .d0(n1667), .sl(n1650), .d1(n1376) );
	nor3i_0 U2730 ( .x(n1729), .a(FREEZE), .b(reg_dst_of_EX_2), .c(reg_dst_of_EX_1) );
	inv_5 U2731 ( .x(n1557), .a(reg_dst_of_EX_1) );
	mux2i_5 U2732 ( .x(reg_dst_of_EX_1), .d0(n560), .sl(reg_dst), .d1(n563) );
	inv_6 U2733 ( .x(n4009), .a(n4452) );
	inv_10 U2734 ( .x(IR_opcode_field[2]), .a(n4009) );
	inv_3 U2735 ( .x(n4011), .a(n3950) );
	mux2_4 U2736 ( .x(n1128), .d0(n1657), .sl(n798), .d1(n4012) );
	inv_4 U2737 ( .x(n4012), .a(N462) );
	nand2i_6 U2738 ( .x(n798), .a(n709), .b(n796) );
	inv_10 U2739 ( .x(IR_opcode_field[0]), .a(n4377) );
	inv_2 U274 ( .x(n1667), .a(N519) );
	buf_16 U2740 ( .x(Imm[10]), .a(N6348) );
	buf_14 U2741 ( .x(reg_out_B[25]), .a(n4455) );
	buf_10 U2742 ( .x(Imm[12]), .a(N6352) );
	buf_10 U2743 ( .x(Imm[31]), .a(N6390) );
	buf_14 U2744 ( .x(Imm[8]), .a(N6344) );
	buf_10 U2745 ( .x(reg_out_B[19]), .a(n4456) );
	and2_4 U2746 ( .x(n4390), .a(n3902), .b(n680) );
	buf_10 U2747 ( .x(reg_out_B[0]), .a(n4458) );
	and2_4 U2748 ( .x(n4394), .a(n3911), .b(n680) );
	and2_4 U2749 ( .x(n4410), .a(n3906), .b(n680) );
	mux2i_1 U275 ( .x(n3905), .d0(n1668), .sl(n1650), .d1(n1349) );
	and2_4 U2750 ( .x(n4434), .a(n3897), .b(n680) );
	and2_4 U2751 ( .x(n4422), .a(n3903), .b(n680) );
	and2_4 U2752 ( .x(n4430), .a(n3895), .b(n680) );
	and2_1 U2753 ( .x(n4388), .a(n3913), .b(n680) );
	and2_1 U2754 ( .x(n4392), .a(n3922), .b(n680) );
	and2_1 U2755 ( .x(n4396), .a(n3893), .b(n681) );
	and2_1 U2756 ( .x(n4398), .a(n3918), .b(n681) );
	and2_1 U2757 ( .x(n4400), .a(n3894), .b(n680) );
	and2_1 U2758 ( .x(n4402), .a(n3907), .b(n680) );
	and2_1 U2759 ( .x(n4404), .a(n3916), .b(n680) );
	inv_2 U276 ( .x(n1668), .a(N518) );
	and2_1 U2760 ( .x(n4406), .a(n3896), .b(n680) );
	and2_1 U2761 ( .x(n4408), .a(n3914), .b(n680) );
	and2_1 U2762 ( .x(n4412), .a(n3912), .b(n680) );
	and2_1 U2763 ( .x(n4414), .a(n3899), .b(n680) );
	and2_1 U2764 ( .x(n4416), .a(n3898), .b(n680) );
	and2_1 U2765 ( .x(n4418), .a(n3917), .b(n680) );
	and2_1 U2766 ( .x(n4420), .a(n3908), .b(n680) );
	and2_1 U2767 ( .x(n4424), .a(n3909), .b(n680) );
	and2_1 U2768 ( .x(n4426), .a(n3904), .b(n680) );
	and2_1 U2769 ( .x(n4428), .a(n3915), .b(n680) );
	mux2i_1 U277 ( .x(n3914), .d0(n1659), .sl(n1650), .d1(n1395) );
	and2_1 U2770 ( .x(n4436), .a(n3901), .b(n681) );
	and2_1 U2771 ( .x(n4438), .a(n3920), .b(n681) );
	and2_1 U2772 ( .x(n4440), .a(n3919), .b(n681) );
	and2_1 U2773 ( .x(n4444), .a(n3921), .b(n681) );
	and2_1 U2774 ( .x(n4446), .a(n3900), .b(n681) );
	and2_1 U2775 ( .x(n4448), .a(n3892), .b(n681) );
	and2_1 U2776 ( .x(n4450), .a(n3891), .b(n680) );
	inv_2 U278 ( .x(n1659), .a(N527) );
	nor2_2 U279 ( .x(n1239), .a(___cell__36997_net129247), .b(n1274) );
	buf_14 U28 ( .x(reg_out_A[20]), .a(n3961) );
	inv_2 U280 ( .x(n1274), .a(N5422) );
	inv_2 U281 ( .x(n1292), .a(N5421) );
	inv_2 U282 ( .x(n1281), .a(N5444) );
	inv_2 U283 ( .x(n1503), .a(N5376) );
	inv_2 U284 ( .x(n1509), .a(N5372) );
	aoi222_1 U285 ( .x(n1022), .a(NPC[25]), .b(n1719), .c(n1732), .d(EPC_25),
		.e(Cause_Reg_25), .f(n1803) );
	inv_2 U286 ( .x(n1507), .a(N6041) );
	inv_2 U287 ( .x(n1506), .a(N5374) );
	oai21_1 U288 ( .x(N6749), .a(n641), .b(___cell__36997_net130580), .c(___cell__36997_net127210) );
	mux2_4 U289 ( .x(n641), .d0(___cell__36997_net129388), .sl(___cell__36997_net129354),
		.d1(___cell__36997_net129389) );
	inv_0 U29 ( .x(n1528), .a(NPC[26]) );
	and2_1 U290 ( .x(n677), .a(n3948), .b(n1515) );
	aoi222_1 U291 ( .x(___cell__36997_net127210), .a(NPC[31]), .b(n1719), .c(n1732),
		.d(EPC_31), .e(Cause_Reg_31), .f(n1803) );
	nor2_1 U292 ( .x(n1120), .a(n1776), .b(n778) );
	inv_5 U293 ( .x(IR_latched_10), .a(n1053) );
	nand2i_2 U294 ( .x(n1054), .a(n4371), .b(n642) );
	nand2i_2 U295 ( .x(n1060), .a(n4370), .b(n1718) );
	nor2_1 U296 ( .x(n1102), .a(n1776), .b(n732) );
	nand2i_2 U297 ( .x(n3811), .a(n1102), .b(n764) );
	nand2i_2 U298 ( .x(n1056), .a(n786), .b(n1718) );
	buf_3 U299 ( .x(n910), .a(n951) );
	and2_5 U3 ( .x(n664), .a(___cell__36997_net130214), .b(N6049) );
	inv_2 U30 ( .x(n750), .a(n3979) );
	mux2i_1 U300 ( .x(n3896), .d0(n1677), .sl(n1650), .d1(n1361) );
	inv_2 U301 ( .x(n1677), .a(N509) );
	nor2_1 U302 ( .x(n1101), .a(n705), .b(n775) );
	nand2i_2 U303 ( .x(n1050), .a(n872), .b(n1718) );
	oai21_1 U306 ( .x(N6742), .a(n1020), .b(n678), .c(n1021) );
	inv_5 U307 ( .x(n1020), .a(n1407) );
	aoi222_1 U308 ( .x(n1021), .a(NPC[24]), .b(n1802), .c(n1732), .d(EPC_24),
		.e(Cause_Reg_24), .f(n1803) );
	oai21_1 U309 ( .x(N6746), .a(n1026), .b(n995), .c(n1027) );
	inv_7 U310 ( .x(n1026), .a(n1355) );
	aoi222_1 U311 ( .x(n1027), .a(NPC[28]), .b(n1802), .c(n1732), .d(EPC_28),
		.e(Cause_Reg_28), .f(n1803) );
	mux2i_1 U312 ( .x(n3916), .d0(n1656), .sl(n1650), .d1(n1657) );
	inv_2 U313 ( .x(n1656), .a(N529) );
	mux2i_1 U314 ( .x(n3907), .d0(n1666), .sl(n1650), .d1(n1304) );
	inv_2 U315 ( .x(n1666), .a(N520) );
	oai21_1 U316 ( .x(N6748), .a(___cell__36997_net126005), .b(n995), .c(n1030) );
	inv_4 U318 ( .x(n1362), .a(N438) );
	aoi222_1 U319 ( .x(n1030), .a(NPC[30]), .b(n1802), .c(n1732), .d(EPC_30),
		.e(Cause_Reg_30), .f(n1803) );
	inv_2 U32 ( .x(n1061), .a(IR_latched_14) );
	buf_3 U320 ( .x(n909), .a(n951) );
	mux2i_1 U321 ( .x(n3894), .d0(n1679), .sl(n1650), .d1(n1357) );
	inv_2 U322 ( .x(n1679), .a(N507) );
	oai21_1 U323 ( .x(N6739), .a(n684), .b(___cell__36997_net130580), .c(n1015) );
	aoi222_1 U324 ( .x(n1015), .a(NPC[21]), .b(n1719), .c(n1732), .d(EPC_21),
		.e(Cause_Reg_21), .f(n1803) );
	inv_2 U325 ( .x(___cell__36997_net130580), .a(n677) );
	aoi222_1 U326 ( .x(n1029), .a(NPC[29]), .b(n1719), .c(n1732), .d(EPC_29),
		.e(Cause_Reg_29), .f(n1803) );
	inv_2 U327 ( .x(n678), .a(n677) );
	inv_4 U328 ( .x(n1342), .a(N439) );
	inv_7 U329 ( .x(n1028), .a(n1341) );
	inv_0 U33 ( .x(n1597), .a(IR_latched_input[10]) );
	oai21_1 U330 ( .x(N6747), .a(n1028), .b(n678), .c(n1029) );
	aoi222_1 U331 ( .x(n1017), .a(NPC[22]), .b(n1802), .c(n1732), .d(EPC_22),
		.e(Cause_Reg_22), .f(n1803) );
	nand2_2 U332 ( .x(n995), .a(n3948), .b(n1515) );
	oai21_1 U333 ( .x(N6740), .a(n1016), .b(n995), .c(n1017) );
	oai21_1 U334 ( .x(N6741), .a(n1018), .b(n1777), .c(n1019) );
	inv_5 U335 ( .x(n1018), .a(n1401) );
	aoi222_1 U336 ( .x(n1019), .a(NPC[23]), .b(n1719), .c(n1732), .d(EPC_23),
		.e(Cause_Reg_23), .f(n1803) );
	oai21_1 U337 ( .x(N6738), .a(n640), .b(n1777), .c(n1013) );
	nand2_2 U338 ( .x(n1777), .a(n3948), .b(n1515) );
	aoi222_1 U339 ( .x(n1013), .a(NPC[20]), .b(n1802), .c(n1732), .d(EPC_20),
		.e(Cause_Reg_20), .f(n1803) );
	inv_2 U34 ( .x(IR_latched_9), .a(n1051) );
	mux2i_1 U340 ( .x(n3919), .d0(n1653), .sl(n1650), .d1(n1387) );
	inv_2 U341 ( .x(n1653), .a(N532) );
	oai21_1 U342 ( .x(N6736), .a(n674), .b(n678), .c(n1011) );
	nand2_2 U343 ( .x(n1082), .a(n1718), .b(IR_opcode_field[1]) );
	mux2i_1 U344 ( .x(n3920), .d0(n1652), .sl(n1650), .d1(n1390) );
	inv_2 U345 ( .x(n1652), .a(N533) );
	aoi221_1 U346 ( .x(n1129), .a(Cause_Reg_6), .b(n1803), .c(n1732), .d(EPC_6),
		.e(n1306) );
	oai21_1 U347 ( .x(N6724), .a(n1128), .b(n678), .c(n1129) );
	oai21_1 U348 ( .x(N6737), .a(n639), .b(n995), .c(n1012) );
	mux2_4 U349 ( .x(n639), .d0(n1382), .sl(___cell__36997_net129354), .d1(n1383) );
	mux2i_2 U35 ( .x(n1053), .d0(current_IR_10), .sl(net149680), .d1(IR_latched_input[10]) );
	aoi222_1 U350 ( .x(n1012), .a(NPC[19]), .b(n1719), .c(n1732), .d(EPC_19),
		.e(Cause_Reg_19), .f(n1803) );
	inv_2 U351 ( .x(n1410), .a(N459) );
	oai21_1 U352 ( .x(N6727), .a(n637), .b(___cell__36997_net130580), .c(n1033) );
	inv_2 U353 ( .x(n1396), .a(N464) );
	mux2_4 U354 ( .x(n636), .d0(n1396), .sl(___cell__36997_net129354), .d1(n1397) );
	inv_5 U355 ( .x(n1001), .a(n1398) );
	oai21_1 U356 ( .x(N6730), .a(n1001), .b(___cell__36997_net130580), .c(n1002) );
	oai21_1 U357 ( .x(N6728), .a(n638), .b(n995), .c(n997) );
	mux2_4 U358 ( .x(n638), .d0(n1391), .sl(___cell__36997_net129354), .d1(n1392) );
	inv_2 U359 ( .x(n1391), .a(N458) );
	inv_4 U36 ( .x(IR_latched_3), .a(n849) );
	nand2_2 U361 ( .x(n1068), .a(n642), .b(IR_opcode_field[0]) );
	inv_2 U362 ( .x(n1386), .a(N465) );
	mux2i_1 U363 ( .x(n3918), .d0(n1654), .sl(n1650), .d1(n1397) );
	or3i_2 U364 ( .x(n681), .a(n744), .b(___cell__36997_net125928), .c(n679) );
	aoi222_1 U365 ( .x(n996), .a(NPC[0]), .b(n1719), .c(n1732), .d(EPC_0),
		.e(Cause_Reg_0), .f(n1803) );
	inv_5 U366 ( .x(n1031), .a(n1393) );
	oai21_1 U367 ( .x(N6726), .a(n1031), .b(n1777), .c(n1032) );
	inv_5 U368 ( .x(n1252), .a(n1388) );
	oai21_1 U369 ( .x(N6720), .a(n1252), .b(n1777), .c(n1253) );
	inv_0 U37 ( .x(n1420), .a(IR_latched_input[3]) );
	nor2_4 U370 ( .x(n1105), .a(n705), .b(n1311) );
	nor2_3 U371 ( .x(n1121), .a(n1776), .b(n696) );
	aoi222_1 U372 ( .x(n1131), .a(NPC[1]), .b(n1802), .c(n1732), .d(EPC_1),
		.e(Cause_Reg_1), .f(n1803) );
	nand2i_2 U373 ( .x(n1064), .a(n829), .b(n1718) );
	nand2i_2 U374 ( .x(n1052), .a(n873), .b(n642) );
	nor2_1 U375 ( .x(n1117), .a(n705), .b(n765) );
	nor2_3 U376 ( .x(n1116), .a(n1776), .b(n701) );
	nor2_3 U377 ( .x(n1115), .a(n705), .b(n762) );
	nand2i_2 U378 ( .x(n1042), .a(n886), .b(n642) );
	inv_2 U379 ( .x(n1041), .a(IR_latched_3) );
	inv_14 U38 ( .x(n737), .a(n865) );
	inv_2 U380 ( .x(n1043), .a(IR_latched_4) );
	mux2i_3 U381 ( .x(IR_latched_4), .d0(n1418), .sl(net149680), .d1(n1419) );
	inv_4 U382 ( .x(counter[0]), .a(n4011) );
	ao21_1 U383 ( .x(n2640), .a(intr_slot), .b(n1092), .c(n1093) );
	nand2i_2 U384 ( .x(n1092), .a(delay_slot), .b(n1739) );
	inv_2 U385 ( .x(n1739), .a(n1267) );
	nand2i_2 U386 ( .x(n1093), .a(n1262), .b(___cell__36997_net126604) );
	oai21_1 U387 ( .x(n1034), .a(___cell__36997_net127190), .b(n1263), .c(CLI) );
	inv_5 U388 ( .x(___cell__36997_net130567), .a(___cell__36997_net126604) );
	mux2i_1 U389 ( .x(n2642), .d0(n627), .sl(___cell__36997_net130125), .d1(n813) );
	inv_0 U39 ( .x(n1040), .a(IR_latched_2) );
	mux2i_1 U390 ( .x(n2652), .d0(n617), .sl(___cell__36997_net130125), .d1(n4371) );
	mux2i_1 U391 ( .x(n2655), .d0(n614), .sl(___cell__36997_net130567), .d1(n4370) );
	mux2i_2 U392 ( .x(n2666), .d0(n603), .sl(___cell__36997_net130567), .d1(n654) );
	mux2i_1 U393 ( .x(n2673), .d0(n596), .sl(___cell__36997_net130567), .d1(n1311) );
	mux2i_1 U394 ( .x(n2674), .d0(n595), .sl(___cell__36997_net130125), .d1(n1553) );
	mux2i_1 U395 ( .x(n2675), .d0(n594), .sl(___cell__36997_net130567), .d1(n1552) );
	mux2i_1 U396 ( .x(n2676), .d0(n1294), .sl(___cell__36997_net130125), .d1(n1551) );
	inv_2 U397 ( .x(n1294), .a(EPC_2) );
	inv_2 U398 ( .x(n1276), .a(EPC_3) );
	mux2i_1 U399 ( .x(n2677), .d0(n1276), .sl(___cell__36997_net130567), .d1(n1550) );
	inv_0 U40 ( .x(n1038), .a(IR_latched_0) );
	mux2i_1 U400 ( .x(n2678), .d0(n577), .sl(___cell__36997_net130125), .d1(n1549) );
	mux2i_1 U401 ( .x(n2679), .d0(n576), .sl(___cell__36997_net130567), .d1(n1548) );
	mux2i_1 U402 ( .x(n2680), .d0(n575), .sl(___cell__36997_net130125), .d1(n1308) );
	mux2i_1 U403 ( .x(n2681), .d0(n574), .sl(___cell__36997_net130567), .d1(n1547) );
	mux2i_1 U404 ( .x(n2682), .d0(n573), .sl(___cell__36997_net130125), .d1(n1546) );
	mux2i_1 U405 ( .x(n2683), .d0(n572), .sl(___cell__36997_net130567), .d1(n1545) );
	mux2i_1 U406 ( .x(n2684), .d0(n593), .sl(___cell__36997_net130125), .d1(n1544) );
	mux2i_1 U407 ( .x(n2685), .d0(n592), .sl(___cell__36997_net130567), .d1(n1543) );
	mux2i_1 U408 ( .x(n2686), .d0(n591), .sl(___cell__36997_net130125), .d1(n1542) );
	mux2i_1 U409 ( .x(n2687), .d0(n590), .sl(___cell__36997_net130567), .d1(n1541) );
	inv_2 U41 ( .x(n824), .a(n1427) );
	mux2i_1 U410 ( .x(n2688), .d0(n589), .sl(___cell__36997_net130125), .d1(n1540) );
	mux2i_1 U411 ( .x(n2689), .d0(n588), .sl(___cell__36997_net130567), .d1(n1539) );
	mux2i_1 U412 ( .x(n2690), .d0(n587), .sl(___cell__36997_net130125), .d1(n1538) );
	mux2i_1 U413 ( .x(n2691), .d0(n586), .sl(___cell__36997_net130567), .d1(n1537) );
	mux2i_1 U414 ( .x(n2692), .d0(n585), .sl(___cell__36997_net130125), .d1(n1536) );
	mux2i_1 U415 ( .x(n2693), .d0(n584), .sl(___cell__36997_net130567), .d1(n1535) );
	mux2i_1 U416 ( .x(n2694), .d0(n583), .sl(___cell__36997_net130567), .d1(n1534) );
	mux2i_1 U417 ( .x(n2695), .d0(n1291), .sl(___cell__36997_net130125), .d1(n1533) );
	inv_2 U418 ( .x(n1291), .a(EPC_21) );
	mux2i_1 U419 ( .x(n2696), .d0(n1289), .sl(___cell__36997_net130567), .d1(n1532) );
	inv_2 U420 ( .x(n1289), .a(EPC_22) );
	mux2i_1 U421 ( .x(n2697), .d0(n1287), .sl(___cell__36997_net130125), .d1(n1531) );
	mux2i_1 U422 ( .x(n2698), .d0(n1285), .sl(___cell__36997_net130567), .d1(n1530) );
	inv_2 U423 ( .x(n1285), .a(EPC_24) );
	mux2i_1 U424 ( .x(n2699), .d0(n1283), .sl(___cell__36997_net130125), .d1(n1529) );
	mux2i_1 U425 ( .x(n2700), .d0(n582), .sl(___cell__36997_net130567), .d1(n1528) );
	mux2i_1 U426 ( .x(n2701), .d0(n581), .sl(___cell__36997_net130125), .d1(n1527) );
	mux2i_1 U427 ( .x(n2702), .d0(n580), .sl(___cell__36997_net130567), .d1(n1526) );
	mux2i_1 U428 ( .x(n2703), .d0(n579), .sl(___cell__36997_net130125), .d1(n1525) );
	mux2i_1 U429 ( .x(n2704), .d0(n662), .sl(___cell__36997_net130125), .d1(n1524) );
	inv_0 U43 ( .x(n805), .a(n879) );
	mux2i_1 U430 ( .x(_EPC_reg_31_net69891), .d0(n578), .sl(___cell__36997_net130567),
		.d1(___cell__36997_net129786) );
	inv_5 U431 ( .x(___cell__36997_net130125), .a(___cell__36997_net126604) );
	nor2i_1 U432 ( .x(n1036), .a(n1260), .b(n1261) );
	mux2_2 U433 ( .x(n2709), .d0(_RegFile_31__0), .sl(n1850), .d1(WB_data[0]) );
	mux2_2 U434 ( .x(n2710), .d0(_RegFile_31__1), .sl(n1850), .d1(WB_data[1]) );
	mux2_2 U435 ( .x(n2711), .d0(_RegFile_31__2), .sl(n1850), .d1(WB_data[2]) );
	mux2_2 U436 ( .x(n2712), .d0(_RegFile_31__3), .sl(n1850), .d1(WB_data[3]) );
	mux2_2 U437 ( .x(n2713), .d0(_RegFile_31__4), .sl(n1850), .d1(WB_data[4]) );
	mux2_2 U438 ( .x(n2714), .d0(_RegFile_31__5), .sl(n1850), .d1(WB_data[5]) );
	mux2_2 U439 ( .x(n2715), .d0(_RegFile_31__6), .sl(n1850), .d1(WB_data[6]) );
	and3_3 U44 ( .x(n1443), .a(n770), .b(n1693), .c(n1692) );
	mux2_2 U440 ( .x(n2716), .d0(_RegFile_31__7), .sl(n1850), .d1(WB_data[7]) );
	mux2i_1 U441 ( .x(n2718), .d0(n2463), .sl(n1850), .d1(n1801) );
	mux2i_1 U442 ( .x(n2719), .d0(n2440), .sl(n1850), .d1(n1778) );
	mux2i_1 U443 ( .x(n2720), .d0(n2441), .sl(n1850), .d1(n1779) );
	mux2i_1 U444 ( .x(n2721), .d0(n2442), .sl(n1850), .d1(n1780) );
	mux2i_1 U445 ( .x(n2722), .d0(n2443), .sl(n1850), .d1(n1781) );
	mux2i_1 U446 ( .x(n2723), .d0(n2444), .sl(n1850), .d1(n1782) );
	mux2i_1 U447 ( .x(n2724), .d0(n2445), .sl(n1850), .d1(n1783) );
	mux2i_1 U448 ( .x(n2725), .d0(n2446), .sl(n1850), .d1(n1784) );
	mux2i_1 U449 ( .x(n2726), .d0(n2447), .sl(n1850), .d1(n1785) );
	mux2i_1 U450 ( .x(n2727), .d0(n2448), .sl(n1850), .d1(n1786) );
	mux2i_1 U451 ( .x(n2728), .d0(n2449), .sl(n1850), .d1(n1787) );
	mux2i_1 U452 ( .x(n2729), .d0(n2450), .sl(n1850), .d1(n1788) );
	mux2i_1 U453 ( .x(n2730), .d0(n2451), .sl(n1850), .d1(n1789) );
	mux2i_1 U454 ( .x(n2731), .d0(n2452), .sl(n1850), .d1(n1790) );
	mux2i_1 U455 ( .x(n2732), .d0(n2453), .sl(n1850), .d1(n1791) );
	mux2i_1 U456 ( .x(n2733), .d0(n2454), .sl(n1850), .d1(n1792) );
	mux2i_1 U457 ( .x(n2734), .d0(n2455), .sl(n1850), .d1(n1793) );
	mux2i_1 U458 ( .x(n2735), .d0(n2456), .sl(n1850), .d1(n1794) );
	mux2i_1 U459 ( .x(n2736), .d0(n2457), .sl(n1850), .d1(n1795) );
	exor2_1 U46 ( .x(n1692), .a(reg_dst_of_EX_0), .b(n884) );
	mux2i_1 U460 ( .x(n2737), .d0(n2458), .sl(n1850), .d1(n1796) );
	mux2i_1 U461 ( .x(n2738), .d0(n2459), .sl(n1850), .d1(n1797) );
	mux2i_1 U462 ( .x(n2739), .d0(n2460), .sl(n1850), .d1(n1798) );
	or2_2 U463 ( .x(n1748), .a(n3940), .b(n3944) );
	mux2_2 U464 ( .x(n2741), .d0(_RegFile_30__0), .sl(n1849), .d1(WB_data[0]) );
	mux2_2 U465 ( .x(n2742), .d0(_RegFile_30__1), .sl(n1849), .d1(WB_data[1]) );
	mux2_2 U466 ( .x(n2743), .d0(_RegFile_30__2), .sl(n1849), .d1(WB_data[2]) );
	mux2_2 U467 ( .x(n2744), .d0(_RegFile_30__3), .sl(n1849), .d1(WB_data[3]) );
	mux2_2 U468 ( .x(n2745), .d0(_RegFile_30__4), .sl(n1849), .d1(WB_data[4]) );
	mux2_2 U469 ( .x(n2746), .d0(_RegFile_30__5), .sl(n1849), .d1(WB_data[5]) );
	exnor2_1 U47 ( .x(n1441), .a(n772), .b(reg_dst_of_EX_3) );
	mux2_2 U470 ( .x(n2747), .d0(_RegFile_30__6), .sl(n1849), .d1(WB_data[6]) );
	mux2_2 U471 ( .x(n2748), .d0(_RegFile_30__7), .sl(n1849), .d1(WB_data[7]) );
	mux2i_1 U472 ( .x(n2750), .d0(n2439), .sl(n1849), .d1(n1801) );
	mux2i_1 U473 ( .x(n2751), .d0(n2416), .sl(n1849), .d1(n1778) );
	mux2i_1 U474 ( .x(n2752), .d0(n2417), .sl(n1849), .d1(n1779) );
	mux2i_1 U475 ( .x(n2753), .d0(n2418), .sl(n1849), .d1(n1780) );
	mux2i_1 U476 ( .x(n2754), .d0(n2419), .sl(n1849), .d1(n1781) );
	mux2i_1 U477 ( .x(n2755), .d0(n2420), .sl(n1849), .d1(n1782) );
	mux2i_1 U478 ( .x(n2756), .d0(n2421), .sl(n1849), .d1(n1783) );
	mux2i_1 U479 ( .x(n2757), .d0(n2422), .sl(n1849), .d1(n1784) );
	inv_2 U48 ( .x(n1584), .a(n1700) );
	mux2i_1 U480 ( .x(n2758), .d0(n2423), .sl(n1849), .d1(n1785) );
	mux2i_1 U481 ( .x(n2759), .d0(n2424), .sl(n1849), .d1(n1786) );
	mux2i_1 U482 ( .x(n2760), .d0(n2425), .sl(n1849), .d1(n1787) );
	mux2i_1 U483 ( .x(n2761), .d0(n2426), .sl(n1849), .d1(n1788) );
	mux2i_1 U484 ( .x(n2762), .d0(n2427), .sl(n1849), .d1(n1789) );
	mux2i_1 U485 ( .x(n2763), .d0(n2428), .sl(n1849), .d1(n1790) );
	mux2i_1 U486 ( .x(n2764), .d0(n2429), .sl(n1849), .d1(n1791) );
	mux2i_1 U487 ( .x(n2765), .d0(n2430), .sl(n1849), .d1(n1792) );
	mux2i_1 U488 ( .x(n2766), .d0(n2431), .sl(n1849), .d1(n1793) );
	mux2i_1 U489 ( .x(n2767), .d0(n2432), .sl(n1849), .d1(n1794) );
	nand2i_0 U49 ( .x(n1583), .a(IR_opcode_field[2]), .b(n4454) );
	mux2i_1 U490 ( .x(n2768), .d0(n2433), .sl(n1849), .d1(n1795) );
	mux2i_1 U491 ( .x(n2769), .d0(n2434), .sl(n1849), .d1(n1796) );
	mux2i_1 U492 ( .x(n2770), .d0(n2435), .sl(n1849), .d1(n1797) );
	mux2i_1 U493 ( .x(n2771), .d0(n2436), .sl(n1849), .d1(n1798) );
	buf_3 U494 ( .x(n928), .a(n987) );
	or2_2 U495 ( .x(n1749), .a(n3940), .b(n3943) );
	mux2_2 U496 ( .x(n2773), .d0(_RegFile_29__0), .sl(n1847), .d1(WB_data[0]) );
	mux2_2 U497 ( .x(n2774), .d0(_RegFile_29__1), .sl(n1847), .d1(WB_data[1]) );
	mux2_2 U498 ( .x(n2775), .d0(_RegFile_29__2), .sl(n1847), .d1(WB_data[2]) );
	mux2_2 U499 ( .x(n2776), .d0(_RegFile_29__3), .sl(n1847), .d1(WB_data[3]) );
	aoi21_1 U50 ( .x(n1582), .a(IR_opcode_field[1]), .b(n1583), .c(n1584) );
	mux2_2 U500 ( .x(n2777), .d0(_RegFile_29__4), .sl(n1847), .d1(WB_data[4]) );
	mux2_2 U501 ( .x(n2778), .d0(_RegFile_29__5), .sl(n1847), .d1(WB_data[5]) );
	mux2_2 U502 ( .x(n2779), .d0(_RegFile_29__6), .sl(n1847), .d1(WB_data[6]) );
	mux2_2 U503 ( .x(n2780), .d0(_RegFile_29__7), .sl(n1847), .d1(WB_data[7]) );
	mux2i_1 U504 ( .x(n2782), .d0(n2391), .sl(n1847), .d1(n1801) );
	mux2i_1 U505 ( .x(n2783), .d0(n2368), .sl(n1847), .d1(n1778) );
	mux2i_1 U506 ( .x(n2784), .d0(n2369), .sl(n1847), .d1(n1779) );
	mux2i_1 U507 ( .x(n2785), .d0(n2370), .sl(n1847), .d1(n1780) );
	mux2i_1 U508 ( .x(n2786), .d0(n2371), .sl(n1847), .d1(n1781) );
	mux2i_1 U509 ( .x(n2787), .d0(n2372), .sl(n1847), .d1(n1782) );
	nand2i_2 U51 ( .x(n1585), .a(n1320), .b(n1586) );
	mux2i_1 U510 ( .x(n2788), .d0(n2373), .sl(n1847), .d1(n1783) );
	mux2i_1 U511 ( .x(n2789), .d0(n2374), .sl(n1847), .d1(n1784) );
	mux2i_1 U512 ( .x(n2790), .d0(n2375), .sl(n1847), .d1(n1785) );
	mux2i_1 U513 ( .x(n2791), .d0(n2376), .sl(n1847), .d1(n1786) );
	mux2i_1 U514 ( .x(n2792), .d0(n2377), .sl(n1847), .d1(n1787) );
	mux2i_1 U515 ( .x(n2793), .d0(n2378), .sl(n1847), .d1(n1788) );
	mux2i_1 U516 ( .x(n2794), .d0(n2379), .sl(n1847), .d1(n1789) );
	mux2i_1 U517 ( .x(n2795), .d0(n2380), .sl(n1847), .d1(n1790) );
	mux2i_1 U518 ( .x(n2796), .d0(n2381), .sl(n1847), .d1(n1791) );
	mux2i_1 U519 ( .x(n2797), .d0(n2382), .sl(n1847), .d1(n1792) );
	nor2i_1 U52 ( .x(n1320), .a(n1321), .b(n1322) );
	mux2i_1 U520 ( .x(n2798), .d0(n2383), .sl(n1847), .d1(n1793) );
	mux2i_1 U521 ( .x(n2799), .d0(n2384), .sl(n1847), .d1(n1794) );
	mux2i_1 U522 ( .x(n2800), .d0(n2385), .sl(n1847), .d1(n1795) );
	mux2i_1 U523 ( .x(n2801), .d0(n2386), .sl(n1847), .d1(n1796) );
	mux2i_1 U524 ( .x(n2802), .d0(n2387), .sl(n1847), .d1(n1797) );
	mux2i_1 U525 ( .x(n2803), .d0(n2388), .sl(n1847), .d1(n1798) );
	or2_2 U526 ( .x(n1751), .a(n3940), .b(n3942) );
	mux2_2 U527 ( .x(n2805), .d0(_RegFile_28__0), .sl(n1846), .d1(WB_data[0]) );
	mux2_2 U528 ( .x(n2806), .d0(_RegFile_28__1), .sl(n1846), .d1(WB_data[1]) );
	mux2_2 U529 ( .x(n2807), .d0(_RegFile_28__2), .sl(n1846), .d1(WB_data[2]) );
	mux2i_1 U53 ( .x(n1586), .d0(n1580), .sl(IR_opcode_field[1]), .d1(n1581) );
	mux2_2 U530 ( .x(n2808), .d0(_RegFile_28__3), .sl(n1846), .d1(WB_data[3]) );
	mux2_2 U531 ( .x(n2809), .d0(_RegFile_28__4), .sl(n1846), .d1(WB_data[4]) );
	mux2_2 U532 ( .x(n2810), .d0(_RegFile_28__5), .sl(n1846), .d1(WB_data[5]) );
	mux2_2 U533 ( .x(n2811), .d0(_RegFile_28__6), .sl(n1846), .d1(WB_data[6]) );
	mux2_2 U534 ( .x(n2812), .d0(_RegFile_28__7), .sl(n1846), .d1(WB_data[7]) );
	mux2i_1 U535 ( .x(n2814), .d0(n2367), .sl(n1846), .d1(n1801) );
	mux2i_1 U536 ( .x(n2815), .d0(n2344), .sl(n1846), .d1(n1778) );
	mux2i_1 U537 ( .x(n2816), .d0(n2345), .sl(n1846), .d1(n1779) );
	mux2i_1 U538 ( .x(n2817), .d0(n2346), .sl(n1846), .d1(n1780) );
	mux2i_1 U539 ( .x(n2818), .d0(n2347), .sl(n1846), .d1(n1781) );
	inv_10 U54 ( .x(___cell__36997_net129477), .a(n331) );
	mux2i_1 U540 ( .x(n2819), .d0(n2348), .sl(n1846), .d1(n1782) );
	mux2i_1 U541 ( .x(n2820), .d0(n2349), .sl(n1846), .d1(n1783) );
	mux2i_1 U542 ( .x(n2821), .d0(n2350), .sl(n1846), .d1(n1784) );
	mux2i_1 U543 ( .x(n2822), .d0(n2351), .sl(n1846), .d1(n1785) );
	mux2i_1 U544 ( .x(n2823), .d0(n2352), .sl(n1846), .d1(n1786) );
	mux2i_1 U545 ( .x(n2824), .d0(n2353), .sl(n1846), .d1(n1787) );
	mux2i_1 U546 ( .x(n2825), .d0(n2354), .sl(n1846), .d1(n1788) );
	mux2i_1 U547 ( .x(n2826), .d0(n2355), .sl(n1846), .d1(n1789) );
	mux2i_1 U548 ( .x(n2827), .d0(n2356), .sl(n1846), .d1(n1790) );
	mux2i_1 U549 ( .x(n2828), .d0(n2357), .sl(n1846), .d1(n1791) );
	exor2_1 U55 ( .x(___cell__36997_net129979), .a(WB_index_0), .b(n879) );
	mux2i_1 U550 ( .x(n2829), .d0(n2358), .sl(n1846), .d1(n1792) );
	mux2i_1 U551 ( .x(n2830), .d0(n2359), .sl(n1846), .d1(n1793) );
	mux2i_1 U552 ( .x(n2831), .d0(n2360), .sl(n1846), .d1(n1794) );
	mux2i_1 U553 ( .x(n2832), .d0(n2361), .sl(n1846), .d1(n1795) );
	mux2i_1 U554 ( .x(n2833), .d0(n2362), .sl(n1846), .d1(n1796) );
	mux2i_1 U555 ( .x(n2834), .d0(n2363), .sl(n1846), .d1(n1797) );
	mux2i_1 U556 ( .x(n2835), .d0(n2364), .sl(n1846), .d1(n1798) );
	buf_3 U557 ( .x(n931), .a(n987) );
	or2_2 U558 ( .x(n1752), .a(n3940), .b(n3941) );
	mux2_2 U559 ( .x(n2837), .d0(_RegFile_27__0), .sl(n1845), .d1(WB_data[0]) );
	buf_3 U56 ( .x(n715), .a(n332) );
	mux2_2 U560 ( .x(n2838), .d0(_RegFile_27__1), .sl(n1845), .d1(WB_data[1]) );
	mux2_2 U561 ( .x(n2839), .d0(_RegFile_27__2), .sl(n1845), .d1(WB_data[2]) );
	mux2_2 U562 ( .x(n2840), .d0(_RegFile_27__3), .sl(n1845), .d1(WB_data[3]) );
	mux2_2 U563 ( .x(n2841), .d0(_RegFile_27__4), .sl(n1845), .d1(WB_data[4]) );
	mux2_2 U564 ( .x(n2842), .d0(_RegFile_27__5), .sl(n1845), .d1(WB_data[5]) );
	mux2_2 U565 ( .x(n2843), .d0(_RegFile_27__6), .sl(n1845), .d1(WB_data[6]) );
	mux2_2 U566 ( .x(n2844), .d0(_RegFile_27__7), .sl(n1845), .d1(WB_data[7]) );
	mux2i_1 U567 ( .x(n2846), .d0(n2343), .sl(n1845), .d1(n1801) );
	mux2i_1 U568 ( .x(n2847), .d0(n2320), .sl(n1845), .d1(n1778) );
	mux2i_1 U569 ( .x(n2848), .d0(n2321), .sl(n1845), .d1(n1779) );
	inv_5 U57 ( .x(___cell__36997_net130306), .a(n709) );
	mux2i_1 U570 ( .x(n2849), .d0(n2322), .sl(n1845), .d1(n1780) );
	mux2i_1 U571 ( .x(n2850), .d0(n2323), .sl(n1845), .d1(n1781) );
	mux2i_1 U572 ( .x(n2851), .d0(n2324), .sl(n1845), .d1(n1782) );
	mux2i_1 U573 ( .x(n2852), .d0(n2325), .sl(n1845), .d1(n1783) );
	mux2i_1 U574 ( .x(n2853), .d0(n2326), .sl(n1845), .d1(n1784) );
	mux2i_1 U575 ( .x(n2854), .d0(n2327), .sl(n1845), .d1(n1785) );
	mux2i_1 U576 ( .x(n2855), .d0(n2328), .sl(n1845), .d1(n1786) );
	mux2i_1 U577 ( .x(n2856), .d0(n2329), .sl(n1845), .d1(n1787) );
	mux2i_1 U578 ( .x(n2857), .d0(n2330), .sl(n1845), .d1(n1788) );
	mux2i_1 U579 ( .x(n2858), .d0(n2331), .sl(n1845), .d1(n1789) );
	mux2i_1 U58 ( .x(n1452), .d0(n628), .sl(opcode_of_MEM_5), .d1(n1579) );
	mux2i_1 U580 ( .x(n2859), .d0(n2332), .sl(n1845), .d1(n1790) );
	mux2i_1 U581 ( .x(n2860), .d0(n2333), .sl(n1845), .d1(n1791) );
	mux2i_1 U582 ( .x(n2861), .d0(n2334), .sl(n1845), .d1(n1792) );
	mux2i_1 U583 ( .x(n2862), .d0(n2335), .sl(n1845), .d1(n1793) );
	mux2i_1 U584 ( .x(n2863), .d0(n2336), .sl(n1845), .d1(n1794) );
	mux2i_1 U585 ( .x(n2864), .d0(n2337), .sl(n1845), .d1(n1795) );
	mux2i_1 U586 ( .x(n2865), .d0(n2338), .sl(n1845), .d1(n1796) );
	mux2i_1 U587 ( .x(n2866), .d0(n2339), .sl(n1845), .d1(n1797) );
	mux2i_1 U588 ( .x(n2867), .d0(n2340), .sl(n1845), .d1(n1798) );
	or2_2 U589 ( .x(n1753), .a(n3939), .b(n3944) );
	nand2i_2 U59 ( .x(n1478), .a(opcode_of_MEM_1), .b(n1690) );
	mux2_2 U590 ( .x(n2869), .d0(_RegFile_26__0), .sl(n1844), .d1(WB_data[0]) );
	mux2_2 U591 ( .x(n2870), .d0(_RegFile_26__1), .sl(n1844), .d1(WB_data[1]) );
	mux2_2 U592 ( .x(n2871), .d0(_RegFile_26__2), .sl(n1844), .d1(WB_data[2]) );
	mux2_2 U593 ( .x(n2872), .d0(_RegFile_26__3), .sl(n1844), .d1(WB_data[3]) );
	mux2_2 U594 ( .x(n2873), .d0(_RegFile_26__4), .sl(n1844), .d1(WB_data[4]) );
	mux2_2 U595 ( .x(n2874), .d0(_RegFile_26__5), .sl(n1844), .d1(WB_data[5]) );
	mux2_2 U596 ( .x(n2875), .d0(_RegFile_26__6), .sl(n1844), .d1(WB_data[6]) );
	mux2_2 U597 ( .x(n2876), .d0(_RegFile_26__7), .sl(n1844), .d1(WB_data[7]) );
	mux2i_1 U598 ( .x(n2878), .d0(n2319), .sl(n1844), .d1(n1801) );
	mux2i_1 U599 ( .x(n2879), .d0(n2296), .sl(n1844), .d1(n1778) );
	inv_2 U60 ( .x(n1690), .a(n1450) );
	mux2i_1 U600 ( .x(n2880), .d0(n2297), .sl(n1844), .d1(n1779) );
	mux2i_1 U601 ( .x(n2881), .d0(n2298), .sl(n1844), .d1(n1780) );
	mux2i_1 U602 ( .x(n2882), .d0(n2299), .sl(n1844), .d1(n1781) );
	mux2i_1 U603 ( .x(n2883), .d0(n2300), .sl(n1844), .d1(n1782) );
	mux2i_1 U604 ( .x(n2884), .d0(n2301), .sl(n1844), .d1(n1783) );
	mux2i_1 U605 ( .x(n2885), .d0(n2302), .sl(n1844), .d1(n1784) );
	mux2i_1 U606 ( .x(n2886), .d0(n2303), .sl(n1844), .d1(n1785) );
	mux2i_1 U607 ( .x(n2887), .d0(n2304), .sl(n1844), .d1(n1786) );
	mux2i_1 U608 ( .x(n2888), .d0(n2305), .sl(n1844), .d1(n1787) );
	mux2i_1 U609 ( .x(n2889), .d0(n2306), .sl(n1844), .d1(n1788) );
	nand2i_2 U61 ( .x(n1450), .a(opcode_of_MEM_5), .b(opcode_of_MEM_3) );
	mux2i_1 U610 ( .x(n2890), .d0(n2307), .sl(n1844), .d1(n1789) );
	mux2i_1 U611 ( .x(n2891), .d0(n2308), .sl(n1844), .d1(n1790) );
	mux2i_1 U612 ( .x(n2892), .d0(n2309), .sl(n1844), .d1(n1791) );
	mux2i_1 U613 ( .x(n2893), .d0(n2310), .sl(n1844), .d1(n1792) );
	mux2i_1 U614 ( .x(n2894), .d0(n2311), .sl(n1844), .d1(n1793) );
	mux2i_1 U615 ( .x(n2895), .d0(n2312), .sl(n1844), .d1(n1794) );
	mux2i_1 U616 ( .x(n2896), .d0(n2313), .sl(n1844), .d1(n1795) );
	mux2i_1 U617 ( .x(n2897), .d0(n2314), .sl(n1844), .d1(n1796) );
	mux2i_1 U618 ( .x(n2898), .d0(n2315), .sl(n1844), .d1(n1797) );
	mux2i_1 U619 ( .x(n2899), .d0(n2316), .sl(n1844), .d1(n1798) );
	and3i_3 U62 ( .x(n1458), .a(n667), .b(n1567), .c(n1566) );
	buf_3 U620 ( .x(n933), .a(n961) );
	or2_2 U621 ( .x(n1754), .a(n3939), .b(n3943) );
	mux2_2 U622 ( .x(n2901), .d0(_RegFile_25__0), .sl(n1843), .d1(WB_data[0]) );
	mux2_2 U623 ( .x(n2902), .d0(_RegFile_25__1), .sl(n1843), .d1(WB_data[1]) );
	mux2_2 U624 ( .x(n2903), .d0(_RegFile_25__2), .sl(n1843), .d1(WB_data[2]) );
	mux2_2 U625 ( .x(n2904), .d0(_RegFile_25__3), .sl(n1843), .d1(WB_data[3]) );
	mux2_2 U626 ( .x(n2905), .d0(_RegFile_25__4), .sl(n1843), .d1(WB_data[4]) );
	mux2_2 U627 ( .x(n2906), .d0(_RegFile_25__5), .sl(n1843), .d1(WB_data[5]) );
	mux2_2 U628 ( .x(n2907), .d0(_RegFile_25__6), .sl(n1843), .d1(WB_data[6]) );
	mux2_2 U629 ( .x(n2908), .d0(_RegFile_25__7), .sl(n1843), .d1(WB_data[7]) );
	exnor2_2 U63 ( .x(n1456), .a(n337), .b(n634) );
	mux2i_1 U630 ( .x(n2910), .d0(n2295), .sl(n1843), .d1(n1801) );
	mux2i_1 U631 ( .x(n2911), .d0(n2272), .sl(n1843), .d1(n1778) );
	mux2i_1 U632 ( .x(n2912), .d0(n2273), .sl(n1843), .d1(n1779) );
	mux2i_1 U633 ( .x(n2913), .d0(n2274), .sl(n1843), .d1(n1780) );
	mux2i_1 U634 ( .x(n2914), .d0(n2275), .sl(n1843), .d1(n1781) );
	mux2i_1 U635 ( .x(n2915), .d0(n2276), .sl(n1843), .d1(n1782) );
	mux2i_1 U636 ( .x(n2916), .d0(n2277), .sl(n1843), .d1(n1783) );
	mux2i_1 U637 ( .x(n2917), .d0(n2278), .sl(n1843), .d1(n1784) );
	mux2i_1 U638 ( .x(n2918), .d0(n2279), .sl(n1843), .d1(n1785) );
	mux2i_1 U639 ( .x(n2919), .d0(n2280), .sl(n1843), .d1(n1786) );
	nand2i_2 U64 ( .x(n1723), .a(n3888), .b(WB_data[7]) );
	mux2i_1 U640 ( .x(n2920), .d0(n2281), .sl(n1843), .d1(n1787) );
	mux2i_1 U641 ( .x(n2921), .d0(n2282), .sl(n1843), .d1(n1788) );
	mux2i_1 U642 ( .x(n2922), .d0(n2283), .sl(n1843), .d1(n1789) );
	mux2i_1 U643 ( .x(n2923), .d0(n2284), .sl(n1843), .d1(n1790) );
	mux2i_1 U644 ( .x(n2924), .d0(n2285), .sl(n1843), .d1(n1791) );
	mux2i_1 U645 ( .x(n2925), .d0(n2286), .sl(n1843), .d1(n1792) );
	mux2i_1 U646 ( .x(n2926), .d0(n2287), .sl(n1843), .d1(n1793) );
	mux2i_1 U647 ( .x(n2927), .d0(n2288), .sl(n1843), .d1(n1794) );
	mux2i_1 U648 ( .x(n2928), .d0(n2289), .sl(n1843), .d1(n1795) );
	mux2i_1 U649 ( .x(n2929), .d0(n2290), .sl(n1843), .d1(n1796) );
	nand2i_2 U65 ( .x(n1305), .a(n3888), .b(N13832) );
	mux2i_1 U650 ( .x(n2930), .d0(n2291), .sl(n1843), .d1(n1797) );
	mux2i_1 U651 ( .x(n2931), .d0(n2292), .sl(n1843), .d1(n1798) );
	or2_2 U652 ( .x(n1755), .a(n3939), .b(n3942) );
	mux2_2 U653 ( .x(n2933), .d0(_RegFile_24__0), .sl(n1842), .d1(WB_data[0]) );
	mux2_2 U654 ( .x(n2934), .d0(_RegFile_24__1), .sl(n1842), .d1(WB_data[1]) );
	mux2_2 U655 ( .x(n2935), .d0(_RegFile_24__2), .sl(n1842), .d1(WB_data[2]) );
	mux2_2 U656 ( .x(n2936), .d0(_RegFile_24__3), .sl(n1842), .d1(WB_data[3]) );
	mux2_2 U657 ( .x(n2937), .d0(_RegFile_24__4), .sl(n1842), .d1(WB_data[4]) );
	mux2_2 U658 ( .x(n2938), .d0(_RegFile_24__5), .sl(n1842), .d1(WB_data[5]) );
	mux2_2 U659 ( .x(n2939), .d0(_RegFile_24__6), .sl(n1842), .d1(WB_data[6]) );
	inv_4 U66 ( .x(n881), .a(n1434) );
	mux2_2 U660 ( .x(n2940), .d0(_RegFile_24__7), .sl(n1842), .d1(WB_data[7]) );
	mux2i_1 U661 ( .x(n2942), .d0(n2271), .sl(n1842), .d1(n1801) );
	mux2i_1 U662 ( .x(n2943), .d0(n2248), .sl(n1842), .d1(n1778) );
	mux2i_1 U663 ( .x(n2944), .d0(n2249), .sl(n1842), .d1(n1779) );
	mux2i_1 U664 ( .x(n2945), .d0(n2250), .sl(n1842), .d1(n1780) );
	mux2i_1 U665 ( .x(n2946), .d0(n2251), .sl(n1842), .d1(n1781) );
	mux2i_1 U666 ( .x(n2947), .d0(n2252), .sl(n1842), .d1(n1782) );
	mux2i_1 U667 ( .x(n2948), .d0(n2253), .sl(n1842), .d1(n1783) );
	mux2i_1 U668 ( .x(n2949), .d0(n2254), .sl(n1842), .d1(n1784) );
	mux2i_1 U669 ( .x(n2950), .d0(n2255), .sl(n1842), .d1(n1785) );
	nand2i_2 U67 ( .x(n1470), .a(n724), .b(n1517) );
	mux2i_1 U670 ( .x(n2951), .d0(n2256), .sl(n1842), .d1(n1786) );
	mux2i_1 U671 ( .x(n2952), .d0(n2257), .sl(n1842), .d1(n1787) );
	mux2i_1 U672 ( .x(n2953), .d0(n2258), .sl(n1842), .d1(n1788) );
	mux2i_1 U673 ( .x(n2954), .d0(n2259), .sl(n1842), .d1(n1789) );
	mux2i_1 U674 ( .x(n2955), .d0(n2260), .sl(n1842), .d1(n1790) );
	mux2i_1 U675 ( .x(n2956), .d0(n2261), .sl(n1842), .d1(n1791) );
	mux2i_1 U676 ( .x(n2957), .d0(n2262), .sl(n1842), .d1(n1792) );
	mux2i_1 U677 ( .x(n2958), .d0(n2263), .sl(n1842), .d1(n1793) );
	mux2i_1 U678 ( .x(n2959), .d0(n2264), .sl(n1842), .d1(n1794) );
	mux2i_1 U679 ( .x(n2960), .d0(n2265), .sl(n1842), .d1(n1795) );
	mux2i_1 U68 ( .x(n1460), .d0(FREEZE), .sl(delay_slot), .d1(n1576) );
	mux2i_1 U680 ( .x(n2961), .d0(n2266), .sl(n1842), .d1(n1796) );
	mux2i_1 U681 ( .x(n2962), .d0(n2267), .sl(n1842), .d1(n1797) );
	mux2i_1 U682 ( .x(n2963), .d0(n2268), .sl(n1842), .d1(n1798) );
	or2_2 U683 ( .x(n1756), .a(n3939), .b(n3941) );
	mux2_2 U684 ( .x(n2965), .d0(_RegFile_23__0), .sl(n1841), .d1(WB_data[0]) );
	mux2_2 U685 ( .x(n2966), .d0(_RegFile_23__1), .sl(n1841), .d1(WB_data[1]) );
	mux2_2 U686 ( .x(n2967), .d0(_RegFile_23__2), .sl(n1841), .d1(n686) );
	mux2_2 U687 ( .x(n2968), .d0(_RegFile_23__3), .sl(n1841), .d1(n685) );
	mux2_2 U688 ( .x(n2969), .d0(_RegFile_23__4), .sl(n1841), .d1(WB_data[4]) );
	mux2_2 U689 ( .x(n2970), .d0(_RegFile_23__5), .sl(n1841), .d1(WB_data[5]) );
	nand2_0 U69 ( .x(n1715), .a(n807), .b(n1462) );
	mux2_2 U690 ( .x(n2971), .d0(_RegFile_23__6), .sl(n1841), .d1(WB_data[6]) );
	mux2_2 U691 ( .x(n2972), .d0(_RegFile_23__7), .sl(n1841), .d1(WB_data[7]) );
	mux2i_1 U692 ( .x(n2974), .d0(n2247), .sl(n1841), .d1(n1801) );
	mux2i_1 U693 ( .x(n2975), .d0(n2224), .sl(n1841), .d1(n1778) );
	mux2i_1 U694 ( .x(n2976), .d0(n2225), .sl(n1841), .d1(n1779) );
	mux2i_1 U695 ( .x(n2977), .d0(n2226), .sl(n1841), .d1(n1780) );
	mux2i_1 U696 ( .x(n2978), .d0(n2227), .sl(n1841), .d1(n1781) );
	mux2i_1 U697 ( .x(n2979), .d0(n2228), .sl(n1841), .d1(n1782) );
	mux2i_1 U698 ( .x(n2980), .d0(n2229), .sl(n1841), .d1(n1783) );
	mux2i_1 U699 ( .x(n2981), .d0(n2230), .sl(n1841), .d1(n1784) );
	mux2i_1 U70 ( .x(n1265), .d0(n1312), .sl(n1454), .d1(n1591) );
	mux2i_1 U700 ( .x(n2982), .d0(n2231), .sl(n1841), .d1(n1785) );
	mux2i_1 U701 ( .x(n2983), .d0(n2232), .sl(n1841), .d1(n1786) );
	mux2i_1 U702 ( .x(n2984), .d0(n2233), .sl(n1841), .d1(n1787) );
	mux2i_1 U703 ( .x(n2985), .d0(n2234), .sl(n1841), .d1(n1788) );
	mux2i_1 U704 ( .x(n2986), .d0(n2235), .sl(n1841), .d1(n1789) );
	mux2i_1 U705 ( .x(n2987), .d0(n2236), .sl(n1841), .d1(n1790) );
	mux2i_1 U706 ( .x(n2988), .d0(n2237), .sl(n1841), .d1(n1791) );
	mux2i_1 U707 ( .x(n2989), .d0(n2238), .sl(n1841), .d1(n1792) );
	mux2i_1 U708 ( .x(n2990), .d0(n2239), .sl(n1841), .d1(n1793) );
	mux2i_1 U709 ( .x(n2991), .d0(n2240), .sl(n1841), .d1(n1794) );
	inv_5 U71 ( .x(n1454), .a(n1440) );
	mux2i_1 U710 ( .x(n2992), .d0(n2241), .sl(n1841), .d1(n1795) );
	mux2i_1 U711 ( .x(n2993), .d0(n2242), .sl(n1841), .d1(n1796) );
	mux2i_1 U712 ( .x(n2994), .d0(n2243), .sl(n1841), .d1(n1797) );
	mux2i_1 U713 ( .x(n2995), .d0(n2244), .sl(n1841), .d1(n1798) );
	or2_2 U714 ( .x(n1757), .a(n3938), .b(n3944) );
	mux2_2 U715 ( .x(n2997), .d0(_RegFile_22__0), .sl(n1840), .d1(WB_data[0]) );
	mux2_2 U716 ( .x(n2998), .d0(_RegFile_22__1), .sl(n1840), .d1(WB_data[1]) );
	mux2_2 U717 ( .x(n2999), .d0(_RegFile_22__2), .sl(n1840), .d1(WB_data[2]) );
	mux2_2 U718 ( .x(n3000), .d0(_RegFile_22__3), .sl(n1840), .d1(WB_data[3]) );
	mux2_2 U719 ( .x(n3001), .d0(_RegFile_22__4), .sl(n1840), .d1(WB_data[4]) );
	nor2_1 U72 ( .x(n1720), .a(n1492), .b(n1484) );
	mux2_2 U720 ( .x(n3002), .d0(_RegFile_22__5), .sl(n1840), .d1(WB_data[5]) );
	mux2_2 U721 ( .x(n3003), .d0(_RegFile_22__6), .sl(n1840), .d1(WB_data[6]) );
	mux2_2 U722 ( .x(n3004), .d0(_RegFile_22__7), .sl(n1840), .d1(WB_data[7]) );
	mux2i_1 U723 ( .x(n3006), .d0(n2223), .sl(n1840), .d1(n1801) );
	mux2i_1 U724 ( .x(n3007), .d0(n2200), .sl(n1840), .d1(n1778) );
	mux2i_1 U725 ( .x(n3008), .d0(n2201), .sl(n1840), .d1(n1779) );
	mux2i_1 U726 ( .x(n3009), .d0(n2202), .sl(n1840), .d1(n1780) );
	mux2i_1 U727 ( .x(n3010), .d0(n2203), .sl(n1840), .d1(n1781) );
	mux2i_1 U728 ( .x(n3011), .d0(n2204), .sl(n1840), .d1(n1782) );
	mux2i_1 U729 ( .x(n3012), .d0(n2205), .sl(n1840), .d1(n1783) );
	nand2i_2 U73 ( .x(n1721), .a(___cell__36997_net125928), .b(n1720) );
	mux2i_1 U730 ( .x(n3013), .d0(n2206), .sl(n1840), .d1(n1784) );
	mux2i_1 U731 ( .x(n3014), .d0(n2207), .sl(n1840), .d1(n1785) );
	mux2i_1 U732 ( .x(n3015), .d0(n2208), .sl(n1840), .d1(n1786) );
	mux2i_1 U733 ( .x(n3016), .d0(n2209), .sl(n1840), .d1(n1787) );
	mux2i_1 U734 ( .x(n3017), .d0(n2210), .sl(n1840), .d1(n1788) );
	mux2i_1 U735 ( .x(n3018), .d0(n2211), .sl(n1840), .d1(n1789) );
	mux2i_1 U736 ( .x(n3019), .d0(n2212), .sl(n1840), .d1(n1790) );
	mux2i_1 U737 ( .x(n3020), .d0(n2213), .sl(n1840), .d1(n1791) );
	mux2i_1 U738 ( .x(n3021), .d0(n2214), .sl(n1840), .d1(n1792) );
	mux2i_1 U739 ( .x(n3022), .d0(n2215), .sl(n1840), .d1(n1793) );
	inv_2 U74 ( .x(n1057), .a(IR_latched_12) );
	mux2i_1 U740 ( .x(n3023), .d0(n2216), .sl(n1840), .d1(n1794) );
	mux2i_1 U741 ( .x(n3024), .d0(n2217), .sl(n1840), .d1(n1795) );
	mux2i_1 U742 ( .x(n3025), .d0(n2218), .sl(n1840), .d1(n1796) );
	mux2i_1 U743 ( .x(n3026), .d0(n2219), .sl(n1840), .d1(n1797) );
	mux2i_1 U744 ( .x(n3027), .d0(n2220), .sl(n1840), .d1(n1798) );
	or2_2 U745 ( .x(n1758), .a(n3938), .b(n3943) );
	mux2_2 U746 ( .x(n3029), .d0(_RegFile_21__0), .sl(n1839), .d1(WB_data[0]) );
	mux2_2 U747 ( .x(n3030), .d0(_RegFile_21__1), .sl(n1839), .d1(WB_data[1]) );
	mux2_2 U748 ( .x(n3031), .d0(_RegFile_21__2), .sl(n1839), .d1(WB_data[2]) );
	mux2_2 U749 ( .x(n3032), .d0(_RegFile_21__3), .sl(n1839), .d1(WB_data[3]) );
	inv_2 U75 ( .x(n1498), .a(N5379) );
	mux2_2 U750 ( .x(n3033), .d0(_RegFile_21__4), .sl(n1839), .d1(WB_data[4]) );
	mux2_2 U751 ( .x(n3034), .d0(_RegFile_21__5), .sl(n1839), .d1(WB_data[5]) );
	mux2_2 U752 ( .x(n3035), .d0(_RegFile_21__6), .sl(n1839), .d1(WB_data[6]) );
	mux2_2 U753 ( .x(n3036), .d0(_RegFile_21__7), .sl(n1839), .d1(WB_data[7]) );
	mux2i_1 U754 ( .x(n3038), .d0(n2199), .sl(n1839), .d1(n1801) );
	mux2i_1 U755 ( .x(n3039), .d0(n2176), .sl(n1839), .d1(n1778) );
	mux2i_1 U756 ( .x(n3040), .d0(n2177), .sl(n1839), .d1(n1779) );
	mux2i_1 U757 ( .x(n3041), .d0(n2178), .sl(n1839), .d1(n1780) );
	mux2i_1 U758 ( .x(n3042), .d0(n2179), .sl(n1839), .d1(n1781) );
	mux2i_1 U759 ( .x(n3043), .d0(n2180), .sl(n1839), .d1(n1782) );
	nand2i_2 U76 ( .x(n1587), .a(n557), .b(n1738) );
	mux2i_1 U760 ( .x(n3044), .d0(n2181), .sl(n1839), .d1(n1783) );
	mux2i_1 U761 ( .x(n3045), .d0(n2182), .sl(n1839), .d1(n1784) );
	mux2i_1 U762 ( .x(n3046), .d0(n2183), .sl(n1839), .d1(n1785) );
	mux2i_1 U763 ( .x(n3047), .d0(n2184), .sl(n1839), .d1(n1786) );
	mux2i_1 U764 ( .x(n3048), .d0(n2185), .sl(n1839), .d1(n1787) );
	mux2i_1 U765 ( .x(n3049), .d0(n2186), .sl(n1839), .d1(n1788) );
	mux2i_1 U766 ( .x(n3050), .d0(n2187), .sl(n1839), .d1(n1789) );
	mux2i_1 U767 ( .x(n3051), .d0(n2188), .sl(n1839), .d1(n1790) );
	mux2i_1 U768 ( .x(n3052), .d0(n2189), .sl(n1839), .d1(n1791) );
	mux2i_1 U769 ( .x(n3053), .d0(n2190), .sl(n1839), .d1(n1792) );
	nand2i_2 U77 ( .x(n1589), .a(___cell__36997_net130681), .b(n1738) );
	mux2i_1 U770 ( .x(n3054), .d0(n2191), .sl(n1839), .d1(n1793) );
	mux2i_1 U771 ( .x(n3055), .d0(n2192), .sl(n1839), .d1(n1794) );
	mux2i_1 U772 ( .x(n3056), .d0(n2193), .sl(n1839), .d1(n1795) );
	mux2i_1 U773 ( .x(n3057), .d0(n2194), .sl(n1839), .d1(n1796) );
	mux2i_1 U774 ( .x(n3058), .d0(n2195), .sl(n1839), .d1(n1797) );
	buf_3 U775 ( .x(n965), .a(n952) );
	mux2i_1 U776 ( .x(n3059), .d0(n2196), .sl(n1839), .d1(n1798) );
	or2_2 U777 ( .x(n1759), .a(n3938), .b(n3942) );
	mux2_2 U778 ( .x(n3061), .d0(_RegFile_20__0), .sl(n1838), .d1(WB_data[0]) );
	mux2_2 U779 ( .x(n3062), .d0(_RegFile_20__1), .sl(n1838), .d1(WB_data[1]) );
	nand2i_2 U78 ( .x(n1588), .a(n557), .b(n1472) );
	mux2_2 U780 ( .x(n3063), .d0(_RegFile_20__2), .sl(n1838), .d1(WB_data[2]) );
	mux2_2 U781 ( .x(n3064), .d0(_RegFile_20__3), .sl(n1838), .d1(WB_data[3]) );
	mux2_2 U782 ( .x(n3065), .d0(_RegFile_20__4), .sl(n1838), .d1(WB_data[4]) );
	mux2_2 U783 ( .x(n3066), .d0(_RegFile_20__5), .sl(n1838), .d1(WB_data[5]) );
	mux2_2 U784 ( .x(n3067), .d0(_RegFile_20__6), .sl(n1838), .d1(WB_data[6]) );
	mux2_2 U785 ( .x(n3068), .d0(_RegFile_20__7), .sl(n1838), .d1(WB_data[7]) );
	mux2i_1 U786 ( .x(n3070), .d0(n2175), .sl(n1838), .d1(n1801) );
	mux2i_1 U787 ( .x(n3071), .d0(n2152), .sl(n1838), .d1(n1778) );
	mux2i_1 U788 ( .x(n3072), .d0(n2153), .sl(n1838), .d1(n1779) );
	mux2i_1 U789 ( .x(n3073), .d0(n2154), .sl(n1838), .d1(n1780) );
	or2_2 U79 ( .x(n1472), .a(intr_slot), .b(delay_slot) );
	mux2i_1 U790 ( .x(n3074), .d0(n2155), .sl(n1838), .d1(n1781) );
	mux2i_1 U791 ( .x(n3075), .d0(n2156), .sl(n1838), .d1(n1782) );
	mux2i_1 U792 ( .x(n3076), .d0(n2157), .sl(n1838), .d1(n1783) );
	mux2i_1 U793 ( .x(n3077), .d0(n2158), .sl(n1838), .d1(n1784) );
	mux2i_1 U794 ( .x(n3078), .d0(n2159), .sl(n1838), .d1(n1785) );
	mux2i_1 U795 ( .x(n3079), .d0(n2160), .sl(n1838), .d1(n1786) );
	mux2i_1 U796 ( .x(n3080), .d0(n2161), .sl(n1838), .d1(n1787) );
	mux2i_1 U797 ( .x(n3081), .d0(n2162), .sl(n1838), .d1(n1788) );
	mux2i_1 U798 ( .x(n3082), .d0(n2163), .sl(n1838), .d1(n1789) );
	mux2i_1 U799 ( .x(n3083), .d0(n2164), .sl(n1838), .d1(n1790) );
	inv_2 U80 ( .x(n1738), .a(n1472) );
	mux2i_1 U800 ( .x(n3084), .d0(n2165), .sl(n1838), .d1(n1791) );
	mux2i_1 U801 ( .x(n3085), .d0(n2166), .sl(n1838), .d1(n1792) );
	mux2i_1 U802 ( .x(n3086), .d0(n2167), .sl(n1838), .d1(n1793) );
	mux2i_1 U803 ( .x(n3087), .d0(n2168), .sl(n1838), .d1(n1794) );
	mux2i_1 U804 ( .x(n3088), .d0(n2169), .sl(n1838), .d1(n1795) );
	mux2i_1 U805 ( .x(n3089), .d0(n2170), .sl(n1838), .d1(n1796) );
	mux2i_1 U806 ( .x(n3090), .d0(n2171), .sl(n1838), .d1(n1797) );
	mux2i_1 U807 ( .x(n3091), .d0(n2172), .sl(n1838), .d1(n1798) );
	or2_2 U808 ( .x(n1760), .a(n3938), .b(n3941) );
	mux2_2 U809 ( .x(n3093), .d0(_RegFile_19__0), .sl(n1836), .d1(WB_data[0]) );
	inv_2 U81 ( .x(n1298), .a(N6035) );
	mux2_2 U810 ( .x(n3094), .d0(_RegFile_19__1), .sl(n1836), .d1(WB_data[1]) );
	mux2_2 U811 ( .x(n3095), .d0(_RegFile_19__2), .sl(n1836), .d1(WB_data[2]) );
	mux2_2 U812 ( .x(n3096), .d0(_RegFile_19__3), .sl(n1836), .d1(WB_data[3]) );
	mux2_2 U813 ( .x(n3097), .d0(_RegFile_19__4), .sl(n1836), .d1(WB_data[4]) );
	mux2_2 U814 ( .x(n3098), .d0(_RegFile_19__5), .sl(n1836), .d1(WB_data[5]) );
	mux2_2 U815 ( .x(n3099), .d0(_RegFile_19__6), .sl(n1836), .d1(WB_data[6]) );
	mux2_2 U816 ( .x(n3100), .d0(_RegFile_19__7), .sl(n1836), .d1(WB_data[7]) );
	mux2i_1 U817 ( .x(n3102), .d0(n2127), .sl(n1836), .d1(n1801) );
	mux2i_1 U818 ( .x(n3103), .d0(n2104), .sl(n1836), .d1(n1778) );
	mux2i_1 U819 ( .x(n3104), .d0(n2105), .sl(n1836), .d1(n1779) );
	nor2_1 U82 ( .x(n1297), .a(___cell__36997_net129239), .b(n1298) );
	mux2i_1 U820 ( .x(n3105), .d0(n2106), .sl(n1836), .d1(n1780) );
	mux2i_1 U821 ( .x(n3106), .d0(n2107), .sl(n1836), .d1(n1781) );
	mux2i_1 U822 ( .x(n3107), .d0(n2108), .sl(n1836), .d1(n1782) );
	mux2i_1 U823 ( .x(n3108), .d0(n2109), .sl(n1836), .d1(n1783) );
	mux2i_1 U824 ( .x(n3109), .d0(n2110), .sl(n1836), .d1(n1784) );
	mux2i_1 U825 ( .x(n3110), .d0(n2111), .sl(n1836), .d1(n1785) );
	mux2i_1 U826 ( .x(n3111), .d0(n2112), .sl(n1836), .d1(n1786) );
	mux2i_1 U827 ( .x(n3112), .d0(n2113), .sl(n1836), .d1(n1787) );
	mux2i_1 U828 ( .x(n3113), .d0(n2114), .sl(n1836), .d1(n1788) );
	mux2i_1 U829 ( .x(n3114), .d0(n2115), .sl(n1836), .d1(n1789) );
	nor2i_1 U83 ( .x(n1301), .a(N6018), .b(___cell__36997_net129239) );
	mux2i_1 U830 ( .x(n3115), .d0(n2116), .sl(n1836), .d1(n1790) );
	mux2i_1 U831 ( .x(n3116), .d0(n2117), .sl(n1836), .d1(n1791) );
	mux2i_1 U832 ( .x(n3117), .d0(n2118), .sl(n1836), .d1(n1792) );
	mux2i_1 U833 ( .x(n3118), .d0(n2119), .sl(n1836), .d1(n1793) );
	mux2i_1 U834 ( .x(n3119), .d0(n2120), .sl(n1836), .d1(n1794) );
	mux2i_1 U835 ( .x(n3120), .d0(n2121), .sl(n1836), .d1(n1795) );
	mux2i_1 U836 ( .x(n3121), .d0(n2122), .sl(n1836), .d1(n1796) );
	mux2i_1 U837 ( .x(n3122), .d0(n2123), .sl(n1836), .d1(n1797) );
	mux2i_1 U838 ( .x(n3123), .d0(n2124), .sl(n1836), .d1(n1798) );
	buf_3 U839 ( .x(n940), .a(n961) );
	inv_2 U84 ( .x(n1508), .a(N5373) );
	or2_2 U840 ( .x(n1762), .a(n3934), .b(n3944) );
	mux2_2 U841 ( .x(n3125), .d0(_RegFile_18__0), .sl(n1835), .d1(WB_data[0]) );
	mux2_2 U842 ( .x(n3126), .d0(_RegFile_18__1), .sl(n1835), .d1(WB_data[1]) );
	mux2_2 U843 ( .x(n3127), .d0(_RegFile_18__2), .sl(n1835), .d1(WB_data[2]) );
	mux2_2 U844 ( .x(n3128), .d0(_RegFile_18__3), .sl(n1835), .d1(WB_data[3]) );
	mux2_2 U845 ( .x(n3129), .d0(_RegFile_18__4), .sl(n1835), .d1(WB_data[4]) );
	mux2_2 U846 ( .x(n3130), .d0(_RegFile_18__5), .sl(n1835), .d1(WB_data[5]) );
	mux2_2 U847 ( .x(n3131), .d0(_RegFile_18__6), .sl(n1835), .d1(WB_data[6]) );
	mux2_2 U848 ( .x(n3132), .d0(_RegFile_18__7), .sl(n1835), .d1(WB_data[7]) );
	mux2i_1 U849 ( .x(n3134), .d0(n2103), .sl(n1835), .d1(n1801) );
	mux2i_1 U850 ( .x(n3135), .d0(n2080), .sl(n1835), .d1(n1778) );
	mux2i_1 U851 ( .x(n3136), .d0(n2081), .sl(n1835), .d1(n1779) );
	mux2i_1 U852 ( .x(n3137), .d0(n2082), .sl(n1835), .d1(n1780) );
	mux2i_1 U853 ( .x(n3138), .d0(n2083), .sl(n1835), .d1(n1781) );
	mux2i_1 U854 ( .x(n3139), .d0(n2084), .sl(n1835), .d1(n1782) );
	mux2i_1 U855 ( .x(n3140), .d0(n2085), .sl(n1835), .d1(n1783) );
	mux2i_1 U856 ( .x(n3141), .d0(n2086), .sl(n1835), .d1(n1784) );
	mux2i_1 U857 ( .x(n3142), .d0(n2087), .sl(n1835), .d1(n1785) );
	mux2i_1 U858 ( .x(n3143), .d0(n2088), .sl(n1835), .d1(n1786) );
	mux2i_1 U859 ( .x(n3144), .d0(n2089), .sl(n1835), .d1(n1787) );
	mux2i_1 U860 ( .x(n3145), .d0(n2090), .sl(n1835), .d1(n1788) );
	mux2i_1 U861 ( .x(n3146), .d0(n2091), .sl(n1835), .d1(n1789) );
	mux2i_1 U862 ( .x(n3147), .d0(n2092), .sl(n1835), .d1(n1790) );
	mux2i_1 U863 ( .x(n3148), .d0(n2093), .sl(n1835), .d1(n1791) );
	mux2i_1 U864 ( .x(n3149), .d0(n2094), .sl(n1835), .d1(n1792) );
	mux2i_1 U865 ( .x(n3150), .d0(n2095), .sl(n1835), .d1(n1793) );
	mux2i_1 U866 ( .x(n3151), .d0(n2096), .sl(n1835), .d1(n1794) );
	mux2i_1 U867 ( .x(n3152), .d0(n2097), .sl(n1835), .d1(n1795) );
	mux2i_1 U868 ( .x(n3153), .d0(n2098), .sl(n1835), .d1(n1796) );
	mux2i_1 U869 ( .x(n3154), .d0(n2099), .sl(n1835), .d1(n1797) );
	mux2i_1 U870 ( .x(n3155), .d0(n2100), .sl(n1835), .d1(n1798) );
	buf_3 U871 ( .x(n941), .a(n961) );
	or2_2 U872 ( .x(n1763), .a(n3934), .b(n3943) );
	mux2_2 U873 ( .x(n3157), .d0(_RegFile_17__0), .sl(n1834), .d1(WB_data[0]) );
	mux2_2 U874 ( .x(n3158), .d0(_RegFile_17__1), .sl(n1834), .d1(WB_data[1]) );
	mux2_2 U875 ( .x(n3159), .d0(_RegFile_17__2), .sl(n1834), .d1(WB_data[2]) );
	mux2_2 U876 ( .x(n3160), .d0(_RegFile_17__3), .sl(n1834), .d1(WB_data[3]) );
	mux2_2 U877 ( .x(n3161), .d0(_RegFile_17__4), .sl(n1834), .d1(WB_data[4]) );
	mux2_2 U878 ( .x(n3162), .d0(_RegFile_17__5), .sl(n1834), .d1(WB_data[5]) );
	mux2_2 U879 ( .x(n3163), .d0(_RegFile_17__6), .sl(n1834), .d1(WB_data[6]) );
	inv_2 U88 ( .x(___cell__36997_net129388), .a(N437) );
	mux2_2 U880 ( .x(n3164), .d0(_RegFile_17__7), .sl(n1834), .d1(WB_data[7]) );
	mux2i_1 U881 ( .x(n3166), .d0(n2079), .sl(n1834), .d1(n1801) );
	mux2i_1 U882 ( .x(n3167), .d0(n2056), .sl(n1834), .d1(n1778) );
	mux2i_1 U883 ( .x(n3168), .d0(n2057), .sl(n1834), .d1(n1779) );
	mux2i_1 U884 ( .x(n3169), .d0(n2058), .sl(n1834), .d1(n1780) );
	mux2i_1 U885 ( .x(n3170), .d0(n2059), .sl(n1834), .d1(n1781) );
	mux2i_1 U886 ( .x(n3171), .d0(n2060), .sl(n1834), .d1(n1782) );
	mux2i_1 U887 ( .x(n3172), .d0(n2061), .sl(n1834), .d1(n1783) );
	mux2i_1 U888 ( .x(n3173), .d0(n2062), .sl(n1834), .d1(n1784) );
	mux2i_1 U889 ( .x(n3174), .d0(n2063), .sl(n1834), .d1(n1785) );
	mux2i_1 U890 ( .x(n3175), .d0(n2064), .sl(n1834), .d1(n1786) );
	mux2i_1 U891 ( .x(n3176), .d0(n2065), .sl(n1834), .d1(n1787) );
	mux2i_1 U892 ( .x(n3177), .d0(n2066), .sl(n1834), .d1(n1788) );
	mux2i_1 U893 ( .x(n3178), .d0(n2067), .sl(n1834), .d1(n1789) );
	mux2i_1 U894 ( .x(n3179), .d0(n2068), .sl(n1834), .d1(n1790) );
	mux2i_1 U895 ( .x(n3180), .d0(n2069), .sl(n1834), .d1(n1791) );
	mux2i_1 U896 ( .x(n3181), .d0(n2070), .sl(n1834), .d1(n1792) );
	mux2i_1 U897 ( .x(n3182), .d0(n2071), .sl(n1834), .d1(n1793) );
	mux2i_1 U898 ( .x(n3183), .d0(n2072), .sl(n1834), .d1(n1794) );
	mux2i_1 U899 ( .x(n3184), .d0(n2073), .sl(n1834), .d1(n1795) );
	nand2i_2 U90 ( .x(n793), .a(n578), .b(n799) );
	mux2i_1 U900 ( .x(n3185), .d0(n2074), .sl(n1834), .d1(n1796) );
	mux2i_1 U901 ( .x(n3186), .d0(n2075), .sl(n1834), .d1(n1797) );
	mux2i_1 U902 ( .x(n3187), .d0(n2076), .sl(n1834), .d1(n1798) );
	buf_3 U903 ( .x(n942), .a(n934) );
	or2_2 U904 ( .x(n1764), .a(n3934), .b(n3942) );
	mux2_2 U905 ( .x(n3189), .d0(_RegFile_16__0), .sl(n1833), .d1(WB_data[0]) );
	mux2_2 U906 ( .x(n3190), .d0(_RegFile_16__1), .sl(n1833), .d1(WB_data[1]) );
	mux2_2 U907 ( .x(n3191), .d0(_RegFile_16__2), .sl(n1833), .d1(WB_data[2]) );
	mux2_2 U908 ( .x(n3192), .d0(_RegFile_16__3), .sl(n1833), .d1(WB_data[3]) );
	mux2_2 U909 ( .x(n3193), .d0(_RegFile_16__4), .sl(n1833), .d1(WB_data[4]) );
	mux2_2 U910 ( .x(n3194), .d0(_RegFile_16__5), .sl(n1833), .d1(WB_data[5]) );
	mux2_2 U911 ( .x(n3195), .d0(_RegFile_16__6), .sl(n1833), .d1(WB_data[6]) );
	mux2_2 U912 ( .x(n3196), .d0(_RegFile_16__7), .sl(n1833), .d1(WB_data[7]) );
	mux2i_1 U913 ( .x(n3198), .d0(n2055), .sl(n1833), .d1(n1801) );
	mux2i_1 U914 ( .x(n3199), .d0(n2032), .sl(n1833), .d1(n1778) );
	mux2i_1 U915 ( .x(n3200), .d0(n2033), .sl(n1833), .d1(n1779) );
	mux2i_1 U916 ( .x(n3201), .d0(n2034), .sl(n1833), .d1(n1780) );
	mux2i_1 U917 ( .x(n3202), .d0(n2035), .sl(n1833), .d1(n1781) );
	mux2i_1 U918 ( .x(n3203), .d0(n2036), .sl(n1833), .d1(n1782) );
	mux2i_1 U919 ( .x(n3204), .d0(n2037), .sl(n1833), .d1(n1783) );
	nor2_1 U92 ( .x(n1259), .a(delay_slot), .b(n2639) );
	mux2i_1 U920 ( .x(n3205), .d0(n2038), .sl(n1833), .d1(n1784) );
	mux2i_1 U921 ( .x(n3206), .d0(n2039), .sl(n1833), .d1(n1785) );
	mux2i_1 U922 ( .x(n3207), .d0(n2040), .sl(n1833), .d1(n1786) );
	mux2i_1 U923 ( .x(n3208), .d0(n2041), .sl(n1833), .d1(n1787) );
	mux2i_1 U924 ( .x(n3209), .d0(n2042), .sl(n1833), .d1(n1788) );
	mux2i_1 U925 ( .x(n3210), .d0(n2043), .sl(n1833), .d1(n1789) );
	mux2i_1 U926 ( .x(n3211), .d0(n2044), .sl(n1833), .d1(n1790) );
	mux2i_1 U927 ( .x(n3212), .d0(n2045), .sl(n1833), .d1(n1791) );
	mux2i_1 U928 ( .x(n3213), .d0(n2046), .sl(n1833), .d1(n1792) );
	mux2i_1 U929 ( .x(n3214), .d0(n2047), .sl(n1833), .d1(n1793) );
	ao21_3 U93 ( .x(n1590), .a(n1448), .b(n861), .c(n755) );
	mux2i_1 U930 ( .x(n3215), .d0(n2048), .sl(n1833), .d1(n1794) );
	mux2i_1 U931 ( .x(n3216), .d0(n2049), .sl(n1833), .d1(n1795) );
	mux2i_1 U932 ( .x(n3217), .d0(n2050), .sl(n1833), .d1(n1796) );
	mux2i_1 U933 ( .x(n3218), .d0(n2051), .sl(n1833), .d1(n1797) );
	mux2i_1 U934 ( .x(n3219), .d0(n2052), .sl(n1833), .d1(n1798) );
	buf_3 U935 ( .x(n943), .a(n934) );
	or2_2 U936 ( .x(n1765), .a(n3934), .b(n3941) );
	mux2_2 U937 ( .x(n3221), .d0(_RegFile_15__0), .sl(n1832), .d1(WB_data[0]) );
	mux2_2 U938 ( .x(n3222), .d0(_RegFile_15__1), .sl(n1832), .d1(WB_data[1]) );
	mux2_2 U939 ( .x(n3223), .d0(_RegFile_15__2), .sl(n1832), .d1(WB_data[2]) );
	inv_4 U94 ( .x(n1356), .a(N440) );
	mux2_2 U940 ( .x(n3224), .d0(_RegFile_15__3), .sl(n1832), .d1(WB_data[3]) );
	mux2_2 U941 ( .x(n3225), .d0(_RegFile_15__4), .sl(n1832), .d1(WB_data[4]) );
	mux2_2 U942 ( .x(n3226), .d0(_RegFile_15__5), .sl(n1832), .d1(WB_data[5]) );
	mux2_2 U943 ( .x(n3227), .d0(_RegFile_15__6), .sl(n1832), .d1(WB_data[6]) );
	mux2_2 U944 ( .x(n3228), .d0(_RegFile_15__7), .sl(n1832), .d1(WB_data[7]) );
	buf_3 U945 ( .x(n960), .a(n985) );
	mux2i_1 U946 ( .x(n3230), .d0(n2031), .sl(n1832), .d1(n1801) );
	mux2i_1 U947 ( .x(n3231), .d0(n2008), .sl(n1832), .d1(n1778) );
	mux2i_1 U948 ( .x(n3232), .d0(n2009), .sl(n1832), .d1(n1779) );
	mux2i_1 U949 ( .x(n3233), .d0(n2010), .sl(n1832), .d1(n1780) );
	inv_2 U95 ( .x(n1402), .a(N445) );
	mux2i_1 U950 ( .x(n3234), .d0(n2011), .sl(n1832), .d1(n1781) );
	mux2i_1 U951 ( .x(n3235), .d0(n2012), .sl(n1832), .d1(n1782) );
	mux2i_1 U952 ( .x(n3236), .d0(n2013), .sl(n1832), .d1(n1783) );
	mux2i_1 U953 ( .x(n3237), .d0(n2014), .sl(n1832), .d1(n1784) );
	mux2i_1 U954 ( .x(n3238), .d0(n2015), .sl(n1832), .d1(n1785) );
	mux2i_1 U955 ( .x(n3239), .d0(n2016), .sl(n1832), .d1(n1786) );
	mux2i_1 U956 ( .x(n3240), .d0(n2017), .sl(n1832), .d1(n1787) );
	mux2i_1 U957 ( .x(n3241), .d0(n2018), .sl(n1832), .d1(n1788) );
	mux2i_1 U958 ( .x(n3242), .d0(n2019), .sl(n1832), .d1(n1789) );
	mux2i_1 U959 ( .x(n3243), .d0(n2020), .sl(n1832), .d1(n1790) );
	inv_2 U96 ( .x(n1380), .a(N448) );
	mux2i_1 U960 ( .x(n3244), .d0(n2021), .sl(n1832), .d1(n1791) );
	mux2i_1 U961 ( .x(n3245), .d0(n2022), .sl(n1832), .d1(n1792) );
	mux2i_1 U962 ( .x(n3246), .d0(n2023), .sl(n1832), .d1(n1793) );
	mux2i_1 U963 ( .x(n3247), .d0(n2024), .sl(n1832), .d1(n1794) );
	mux2i_1 U964 ( .x(n3248), .d0(n2025), .sl(n1832), .d1(n1795) );
	mux2i_1 U965 ( .x(n3249), .d0(n2026), .sl(n1832), .d1(n1796) );
	mux2i_1 U966 ( .x(n3250), .d0(n2027), .sl(n1832), .d1(n1797) );
	mux2i_1 U967 ( .x(n3251), .d0(n2028), .sl(n1832), .d1(n1798) );
	buf_3 U968 ( .x(n944), .a(n934) );
	or2_2 U969 ( .x(n1766), .a(n3937), .b(n3940) );
	inv_5 U97 ( .x(n1719), .a(n1307) );
	mux2_2 U970 ( .x(n3253), .d0(_RegFile_14__0), .sl(n1831), .d1(WB_data[0]) );
	mux2_2 U971 ( .x(n3254), .d0(_RegFile_14__1), .sl(n1831), .d1(WB_data[1]) );
	mux2_2 U972 ( .x(n3255), .d0(_RegFile_14__2), .sl(n1831), .d1(WB_data[2]) );
	mux2_2 U973 ( .x(n3256), .d0(_RegFile_14__3), .sl(n1831), .d1(WB_data[3]) );
	mux2_2 U974 ( .x(n3257), .d0(_RegFile_14__4), .sl(n1831), .d1(WB_data[4]) );
	mux2_2 U975 ( .x(n3258), .d0(_RegFile_14__5), .sl(n1831), .d1(WB_data[5]) );
	mux2_2 U976 ( .x(n3259), .d0(_RegFile_14__6), .sl(n1831), .d1(WB_data[6]) );
	mux2_2 U977 ( .x(n3260), .d0(_RegFile_14__7), .sl(n1831), .d1(WB_data[7]) );
	mux2i_1 U978 ( .x(n3262), .d0(n2007), .sl(n1831), .d1(n1801) );
	mux2i_1 U979 ( .x(n3263), .d0(n1984), .sl(n1831), .d1(n1778) );
	nand2_1 U98 ( .x(n1307), .a(n1468), .b(___cell__36997_net126612) );
	mux2i_1 U980 ( .x(n3264), .d0(n1985), .sl(n1831), .d1(n1779) );
	mux2i_1 U981 ( .x(n3265), .d0(n1986), .sl(n1831), .d1(n1780) );
	mux2i_1 U982 ( .x(n3266), .d0(n1987), .sl(n1831), .d1(n1781) );
	mux2i_1 U983 ( .x(n3267), .d0(n1988), .sl(n1831), .d1(n1782) );
	mux2i_1 U984 ( .x(n3268), .d0(n1989), .sl(n1831), .d1(n1783) );
	mux2i_1 U985 ( .x(n3269), .d0(n1990), .sl(n1831), .d1(n1784) );
	mux2i_1 U986 ( .x(n3270), .d0(n1991), .sl(n1831), .d1(n1785) );
	mux2i_1 U987 ( .x(n3271), .d0(n1992), .sl(n1831), .d1(n1786) );
	mux2i_1 U988 ( .x(n3272), .d0(n1993), .sl(n1831), .d1(n1787) );
	mux2i_1 U989 ( .x(n3273), .d0(n1994), .sl(n1831), .d1(n1788) );
	nor2_1 U99 ( .x(n1306), .a(n1307), .b(n1308) );
	mux2i_1 U990 ( .x(n3274), .d0(n1995), .sl(n1831), .d1(n1789) );
	mux2i_1 U991 ( .x(n3275), .d0(n1996), .sl(n1831), .d1(n1790) );
	mux2i_1 U992 ( .x(n3276), .d0(n1997), .sl(n1831), .d1(n1791) );
	mux2i_1 U993 ( .x(n3277), .d0(n1998), .sl(n1831), .d1(n1792) );
	mux2i_1 U994 ( .x(n3278), .d0(n1999), .sl(n1831), .d1(n1793) );
	mux2i_1 U995 ( .x(n3279), .d0(n2000), .sl(n1831), .d1(n1794) );
	mux2i_1 U996 ( .x(n3280), .d0(n2001), .sl(n1831), .d1(n1795) );
	mux2i_1 U997 ( .x(n3281), .d0(n2002), .sl(n1831), .d1(n1796) );
	mux2i_1 U998 ( .x(n3282), .d0(n2003), .sl(n1831), .d1(n1797) );
	mux2i_1 U999 ( .x(n3283), .d0(n2004), .sl(n1831), .d1(n1798) );
	smlatnr_1 WB_index_reg_0__master ( .q(WB_index_reg_0__m2s), .qb(), .d(reg_dst_of_MEM_0),
		.sdi(n2461), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 WB_index_reg_0__slave ( .q(WB_index_0), .qb(n3928), .d(WB_index_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 WB_index_reg_1__master ( .q(WB_index_reg_1__m2s), .qb(), .d(reg_dst_of_MEM_1),
		.sdi(n3928), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 WB_index_reg_1__slave ( .q(WB_index_1), .qb(n3929), .d(WB_index_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 WB_index_reg_2__master ( .q(WB_index_reg_2__m2s), .qb(), .d(reg_dst_of_MEM_2),
		.sdi(n3929), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 WB_index_reg_2__slave ( .q(WB_index_2), .qb(n3925), .d(WB_index_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 WB_index_reg_3__master ( .q(WB_index_reg_3__m2s), .qb(), .d(reg_dst_of_MEM_3),
		.sdi(n3925), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 WB_index_reg_3__slave ( .q(WB_index_3), .qb(n3926), .d(WB_index_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 WB_index_reg_4__master ( .q(WB_index_reg_4__m2s), .qb(), .d(reg_dst_of_MEM_4),
		.sdi(WB_index_3), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n913), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 WB_index_reg_4__slave ( .q(WB_index_4), .qb(___cell__6171_net27367),
		.d(WB_index_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__0__master ( .q(_RegFile_reg_0__0__m2s), .qb(),
		.d(n3701), .sdi(n4369), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__0__slave ( .q(_RegFile_0__0), .qb(n4368), .d(_RegFile_reg_0__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__10__master ( .q(_RegFile_reg_0__10__m2s), .qb(),
		.d(n3711), .sdi(n1887), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__10__slave ( .q(_RegFile_0__10), .qb(n1864), .d(_RegFile_reg_0__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__11__master ( .q(_RegFile_reg_0__11__m2s), .qb(),
		.d(n3712), .sdi(n1864), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__11__slave ( .q(_RegFile_0__11), .qb(n1865), .d(_RegFile_reg_0__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__12__master ( .q(_RegFile_reg_0__12__m2s), .qb(),
		.d(n3713), .sdi(n1865), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__12__slave ( .q(_RegFile_0__12), .qb(n1866), .d(_RegFile_reg_0__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__13__master ( .q(_RegFile_reg_0__13__m2s), .qb(),
		.d(n3714), .sdi(n1866), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__13__slave ( .q(_RegFile_0__13), .qb(n1867), .d(_RegFile_reg_0__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__14__master ( .q(_RegFile_reg_0__14__m2s), .qb(),
		.d(n3715), .sdi(n1867), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n955),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__14__slave ( .q(_RegFile_0__14), .qb(n1868), .d(_RegFile_reg_0__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n955), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__15__master ( .q(_RegFile_reg_0__15__m2s), .qb(),
		.d(n3716), .sdi(n1868), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__15__slave ( .q(_RegFile_0__15), .qb(n1869), .d(_RegFile_reg_0__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__16__master ( .q(_RegFile_reg_0__16__m2s), .qb(),
		.d(n3717), .sdi(n1869), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__16__slave ( .q(_RegFile_0__16), .qb(n1870), .d(_RegFile_reg_0__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__17__master ( .q(_RegFile_reg_0__17__m2s), .qb(),
		.d(n3718), .sdi(n1870), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__17__slave ( .q(_RegFile_0__17), .qb(n1871), .d(_RegFile_reg_0__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__18__master ( .q(_RegFile_reg_0__18__m2s), .qb(),
		.d(n3719), .sdi(n1871), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__18__slave ( .q(_RegFile_0__18), .qb(n1872), .d(_RegFile_reg_0__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__19__master ( .q(_RegFile_reg_0__19__m2s), .qb(),
		.d(n3720), .sdi(n1872), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__19__slave ( .q(_RegFile_0__19), .qb(n1873), .d(_RegFile_reg_0__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__1__master ( .q(_RegFile_reg_0__1__m2s), .qb(),
		.d(n3702), .sdi(n4368), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__1__slave ( .q(_RegFile_0__1), .qb(n4367), .d(_RegFile_reg_0__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__20__master ( .q(_RegFile_reg_0__20__m2s), .qb(),
		.d(n3721), .sdi(n1873), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__20__slave ( .q(_RegFile_0__20), .qb(n1874), .d(_RegFile_reg_0__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__21__master ( .q(_RegFile_reg_0__21__m2s), .qb(),
		.d(n3722), .sdi(n1874), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__21__slave ( .q(_RegFile_0__21), .qb(n1875), .d(_RegFile_reg_0__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__22__master ( .q(_RegFile_reg_0__22__m2s), .qb(),
		.d(n3723), .sdi(n1875), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__22__slave ( .q(_RegFile_0__22), .qb(n1876), .d(_RegFile_reg_0__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__23__master ( .q(_RegFile_reg_0__23__m2s), .qb(),
		.d(n3724), .sdi(n1876), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__23__slave ( .q(_RegFile_0__23), .qb(n1877), .d(_RegFile_reg_0__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__24__master ( .q(_RegFile_reg_0__24__m2s), .qb(),
		.d(n3725), .sdi(n1877), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__24__slave ( .q(_RegFile_0__24), .qb(n1878), .d(_RegFile_reg_0__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__25__master ( .q(_RegFile_reg_0__25__m2s), .qb(),
		.d(n3726), .sdi(n1878), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__25__slave ( .q(_RegFile_0__25), .qb(n1879), .d(_RegFile_reg_0__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__26__master ( .q(_RegFile_reg_0__26__m2s), .qb(),
		.d(n3727), .sdi(n1879), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__26__slave ( .q(_RegFile_0__26), .qb(n1880), .d(_RegFile_reg_0__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__27__master ( .q(_RegFile_reg_0__27__m2s), .qb(),
		.d(n3728), .sdi(n1880), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__27__slave ( .q(_RegFile_0__27), .qb(n1881), .d(_RegFile_reg_0__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__28__master ( .q(_RegFile_reg_0__28__m2s), .qb(),
		.d(n3729), .sdi(n1881), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__28__slave ( .q(_RegFile_0__28), .qb(n1882), .d(_RegFile_reg_0__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__29__master ( .q(_RegFile_reg_0__29__m2s), .qb(),
		.d(n3730), .sdi(n1882), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__29__slave ( .q(_RegFile_0__29), .qb(n1883), .d(_RegFile_reg_0__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__2__master ( .q(_RegFile_reg_0__2__m2s), .qb(),
		.d(n3703), .sdi(n4367), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__2__slave ( .q(_RegFile_0__2), .qb(n4366), .d(_RegFile_reg_0__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__30__master ( .q(_RegFile_reg_0__30__m2s), .qb(),
		.d(n3731), .sdi(n1883), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__30__slave ( .q(_RegFile_0__30), .qb(n1884), .d(_RegFile_reg_0__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__31__master ( .q(_RegFile_reg_0__31__m2s), .qb(),
		.d(n3732), .sdi(n1884), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__31__slave ( .q(_RegFile_0__31), .qb(n1885), .d(_RegFile_reg_0__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__3__master ( .q(_RegFile_reg_0__3__m2s), .qb(),
		.d(n3704), .sdi(n4366), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__3__slave ( .q(_RegFile_0__3), .qb(n4365), .d(_RegFile_reg_0__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__4__master ( .q(_RegFile_reg_0__4__m2s), .qb(),
		.d(n3705), .sdi(n4365), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__4__slave ( .q(_RegFile_0__4), .qb(n4364), .d(_RegFile_reg_0__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__5__master ( .q(_RegFile_reg_0__5__m2s), .qb(),
		.d(n3706), .sdi(n4364), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__5__slave ( .q(_RegFile_0__5), .qb(n4363), .d(_RegFile_reg_0__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__6__master ( .q(_RegFile_reg_0__6__m2s), .qb(),
		.d(n3707), .sdi(n4363), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__6__slave ( .q(_RegFile_0__6), .qb(n4362), .d(_RegFile_reg_0__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__7__master ( .q(_RegFile_reg_0__7__m2s), .qb(),
		.d(n3708), .sdi(n4362), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__7__slave ( .q(_RegFile_0__7), .qb(n4361), .d(_RegFile_reg_0__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__8__master ( .q(_RegFile_reg_0__8__m2s), .qb(),
		.d(n3709), .sdi(n4361), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__8__slave ( .q(_RegFile_0__8), .qb(n1886), .d(_RegFile_reg_0__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_0__9__master ( .q(_RegFile_reg_0__9__m2s), .qb(),
		.d(n3710), .sdi(n1886), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_0__9__slave ( .q(_RegFile_0__9), .qb(n1887), .d(_RegFile_reg_0__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__0__master ( .q(_RegFile_reg_10__0__m2s), .qb(),
		.d(n3381), .sdi(n2629), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__0__slave ( .q(_RegFile_10__0), .qb(n4288), .d(_RegFile_reg_10__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__10__master ( .q(_RegFile_reg_10__10__m2s), .qb(),
		.d(n3391), .sdi(n1911), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__10__slave ( .q(_RegFile_10__10), .qb(n1888),
		.d(_RegFile_reg_10__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__11__master ( .q(_RegFile_reg_10__11__m2s), .qb(),
		.d(n3392), .sdi(n1888), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__11__slave ( .q(_RegFile_10__11), .qb(n1889),
		.d(_RegFile_reg_10__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__12__master ( .q(_RegFile_reg_10__12__m2s), .qb(),
		.d(n3393), .sdi(n1889), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n956),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__12__slave ( .q(_RegFile_10__12), .qb(n1890),
		.d(_RegFile_reg_10__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n956), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__13__master ( .q(_RegFile_reg_10__13__m2s), .qb(),
		.d(n3394), .sdi(n1890), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__13__slave ( .q(_RegFile_10__13), .qb(n1891),
		.d(_RegFile_reg_10__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__14__master ( .q(_RegFile_reg_10__14__m2s), .qb(),
		.d(n3395), .sdi(n1891), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__14__slave ( .q(_RegFile_10__14), .qb(n1892),
		.d(_RegFile_reg_10__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__15__master ( .q(_RegFile_reg_10__15__m2s), .qb(),
		.d(n3396), .sdi(n1892), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__15__slave ( .q(_RegFile_10__15), .qb(n1893),
		.d(_RegFile_reg_10__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__16__master ( .q(_RegFile_reg_10__16__m2s), .qb(),
		.d(n3397), .sdi(n1893), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__16__slave ( .q(_RegFile_10__16), .qb(n1894),
		.d(_RegFile_reg_10__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__17__master ( .q(_RegFile_reg_10__17__m2s), .qb(),
		.d(n3398), .sdi(n1894), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__17__slave ( .q(_RegFile_10__17), .qb(n1895),
		.d(_RegFile_reg_10__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__18__master ( .q(_RegFile_reg_10__18__m2s), .qb(),
		.d(n3399), .sdi(n1895), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__18__slave ( .q(_RegFile_10__18), .qb(n1896),
		.d(_RegFile_reg_10__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__19__master ( .q(_RegFile_reg_10__19__m2s), .qb(),
		.d(n3400), .sdi(n1896), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__19__slave ( .q(_RegFile_10__19), .qb(n1897),
		.d(_RegFile_reg_10__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__1__master ( .q(_RegFile_reg_10__1__m2s), .qb(),
		.d(n3382), .sdi(n4288), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__1__slave ( .q(_RegFile_10__1), .qb(n4287), .d(_RegFile_reg_10__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__20__master ( .q(_RegFile_reg_10__20__m2s), .qb(),
		.d(n3401), .sdi(n1897), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__20__slave ( .q(_RegFile_10__20), .qb(n1898),
		.d(_RegFile_reg_10__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__21__master ( .q(_RegFile_reg_10__21__m2s), .qb(),
		.d(n3402), .sdi(n1898), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__21__slave ( .q(_RegFile_10__21), .qb(n1899),
		.d(_RegFile_reg_10__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__22__master ( .q(_RegFile_reg_10__22__m2s), .qb(),
		.d(n3403), .sdi(n1899), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__22__slave ( .q(_RegFile_10__22), .qb(n1900),
		.d(_RegFile_reg_10__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__23__master ( .q(_RegFile_reg_10__23__m2s), .qb(),
		.d(n3404), .sdi(n1900), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__23__slave ( .q(_RegFile_10__23), .qb(n1901),
		.d(_RegFile_reg_10__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__24__master ( .q(_RegFile_reg_10__24__m2s), .qb(),
		.d(n3405), .sdi(n1901), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__24__slave ( .q(_RegFile_10__24), .qb(n1902),
		.d(_RegFile_reg_10__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__25__master ( .q(_RegFile_reg_10__25__m2s), .qb(),
		.d(n3406), .sdi(n1902), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__25__slave ( .q(_RegFile_10__25), .qb(n1903),
		.d(_RegFile_reg_10__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__26__master ( .q(_RegFile_reg_10__26__m2s), .qb(),
		.d(n3407), .sdi(n1903), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__26__slave ( .q(_RegFile_10__26), .qb(n1904),
		.d(_RegFile_reg_10__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__27__master ( .q(_RegFile_reg_10__27__m2s), .qb(),
		.d(n3408), .sdi(n1904), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__27__slave ( .q(_RegFile_10__27), .qb(n1905),
		.d(_RegFile_reg_10__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__28__master ( .q(_RegFile_reg_10__28__m2s), .qb(),
		.d(n3409), .sdi(n1905), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__28__slave ( .q(_RegFile_10__28), .qb(n1906),
		.d(_RegFile_reg_10__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__29__master ( .q(_RegFile_reg_10__29__m2s), .qb(),
		.d(n3410), .sdi(n1906), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__29__slave ( .q(_RegFile_10__29), .qb(n1907),
		.d(_RegFile_reg_10__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__2__master ( .q(_RegFile_reg_10__2__m2s), .qb(),
		.d(n3383), .sdi(n4287), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__2__slave ( .q(_RegFile_10__2), .qb(n4286), .d(_RegFile_reg_10__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__30__master ( .q(_RegFile_reg_10__30__m2s), .qb(),
		.d(n3411), .sdi(n1907), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__30__slave ( .q(_RegFile_10__30), .qb(n1908),
		.d(_RegFile_reg_10__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__31__master ( .q(_RegFile_reg_10__31__m2s), .qb(),
		.d(n3412), .sdi(n1908), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__31__slave ( .q(_RegFile_10__31), .qb(n1909),
		.d(_RegFile_reg_10__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__3__master ( .q(_RegFile_reg_10__3__m2s), .qb(),
		.d(n3384), .sdi(n4286), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__3__slave ( .q(_RegFile_10__3), .qb(n4285), .d(_RegFile_reg_10__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__4__master ( .q(_RegFile_reg_10__4__m2s), .qb(),
		.d(n3385), .sdi(n4285), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__4__slave ( .q(_RegFile_10__4), .qb(n4284), .d(_RegFile_reg_10__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__5__master ( .q(_RegFile_reg_10__5__m2s), .qb(),
		.d(n3386), .sdi(n4284), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__5__slave ( .q(_RegFile_10__5), .qb(n4283), .d(_RegFile_reg_10__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__6__master ( .q(_RegFile_reg_10__6__m2s), .qb(),
		.d(n3387), .sdi(n4283), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__6__slave ( .q(_RegFile_10__6), .qb(n4282), .d(_RegFile_reg_10__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__7__master ( .q(_RegFile_reg_10__7__m2s), .qb(),
		.d(n3388), .sdi(n4282), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__7__slave ( .q(_RegFile_10__7), .qb(n4281), .d(_RegFile_reg_10__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__8__master ( .q(_RegFile_reg_10__8__m2s), .qb(),
		.d(n3389), .sdi(n4281), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__8__slave ( .q(_RegFile_10__8), .qb(n1910), .d(_RegFile_reg_10__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_10__9__master ( .q(_RegFile_reg_10__9__m2s), .qb(),
		.d(n3390), .sdi(n1910), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_10__9__slave ( .q(_RegFile_10__9), .qb(n1911), .d(_RegFile_reg_10__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__0__master ( .q(_RegFile_reg_11__0__m2s), .qb(),
		.d(n3349), .sdi(n1909), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__0__slave ( .q(_RegFile_11__0), .qb(n4280), .d(_RegFile_reg_11__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__10__master ( .q(_RegFile_reg_11__10__m2s), .qb(),
		.d(n3359), .sdi(n1935), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n957),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__10__slave ( .q(_RegFile_11__10), .qb(n1912),
		.d(_RegFile_reg_11__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n957), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__11__master ( .q(_RegFile_reg_11__11__m2s), .qb(),
		.d(n3360), .sdi(n1912), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__11__slave ( .q(_RegFile_11__11), .qb(n1913),
		.d(_RegFile_reg_11__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__12__master ( .q(_RegFile_reg_11__12__m2s), .qb(),
		.d(n3361), .sdi(n1913), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__12__slave ( .q(_RegFile_11__12), .qb(n1914),
		.d(_RegFile_reg_11__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__13__master ( .q(_RegFile_reg_11__13__m2s), .qb(),
		.d(n3362), .sdi(n1914), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__13__slave ( .q(_RegFile_11__13), .qb(n1915),
		.d(_RegFile_reg_11__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__14__master ( .q(_RegFile_reg_11__14__m2s), .qb(),
		.d(n3363), .sdi(n1915), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__14__slave ( .q(_RegFile_11__14), .qb(n1916),
		.d(_RegFile_reg_11__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__15__master ( .q(_RegFile_reg_11__15__m2s), .qb(),
		.d(n3364), .sdi(n1916), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__15__slave ( .q(_RegFile_11__15), .qb(n1917),
		.d(_RegFile_reg_11__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__16__master ( .q(_RegFile_reg_11__16__m2s), .qb(),
		.d(n3365), .sdi(n1917), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__16__slave ( .q(_RegFile_11__16), .qb(n1918),
		.d(_RegFile_reg_11__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__17__master ( .q(_RegFile_reg_11__17__m2s), .qb(),
		.d(n3366), .sdi(n1918), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__17__slave ( .q(_RegFile_11__17), .qb(n1919),
		.d(_RegFile_reg_11__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__18__master ( .q(_RegFile_reg_11__18__m2s), .qb(),
		.d(n3367), .sdi(n1919), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__18__slave ( .q(_RegFile_11__18), .qb(n1920),
		.d(_RegFile_reg_11__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__19__master ( .q(_RegFile_reg_11__19__m2s), .qb(),
		.d(n3368), .sdi(n1920), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__19__slave ( .q(_RegFile_11__19), .qb(n1921),
		.d(_RegFile_reg_11__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__1__master ( .q(_RegFile_reg_11__1__m2s), .qb(),
		.d(n3350), .sdi(n4280), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__1__slave ( .q(_RegFile_11__1), .qb(n4279), .d(_RegFile_reg_11__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__20__master ( .q(_RegFile_reg_11__20__m2s), .qb(),
		.d(n3369), .sdi(n1921), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__20__slave ( .q(_RegFile_11__20), .qb(n1922),
		.d(_RegFile_reg_11__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__21__master ( .q(_RegFile_reg_11__21__m2s), .qb(),
		.d(n3370), .sdi(n1922), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__21__slave ( .q(_RegFile_11__21), .qb(n1923),
		.d(_RegFile_reg_11__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__22__master ( .q(_RegFile_reg_11__22__m2s), .qb(),
		.d(n3371), .sdi(n1923), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__22__slave ( .q(_RegFile_11__22), .qb(n1924),
		.d(_RegFile_reg_11__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__23__master ( .q(_RegFile_reg_11__23__m2s), .qb(),
		.d(n3372), .sdi(n1924), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__23__slave ( .q(_RegFile_11__23), .qb(n1925),
		.d(_RegFile_reg_11__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__24__master ( .q(_RegFile_reg_11__24__m2s), .qb(),
		.d(n3373), .sdi(n1925), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__24__slave ( .q(_RegFile_11__24), .qb(n1926),
		.d(_RegFile_reg_11__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__25__master ( .q(_RegFile_reg_11__25__m2s), .qb(),
		.d(n3374), .sdi(n1926), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__25__slave ( .q(_RegFile_11__25), .qb(n1927),
		.d(_RegFile_reg_11__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__26__master ( .q(_RegFile_reg_11__26__m2s), .qb(),
		.d(n3375), .sdi(n1927), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__26__slave ( .q(_RegFile_11__26), .qb(n1928),
		.d(_RegFile_reg_11__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__27__master ( .q(_RegFile_reg_11__27__m2s), .qb(),
		.d(n3376), .sdi(n1928), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__27__slave ( .q(_RegFile_11__27), .qb(n1929),
		.d(_RegFile_reg_11__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__28__master ( .q(_RegFile_reg_11__28__m2s), .qb(),
		.d(n3377), .sdi(n1929), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__28__slave ( .q(_RegFile_11__28), .qb(n1930),
		.d(_RegFile_reg_11__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__29__master ( .q(_RegFile_reg_11__29__m2s), .qb(),
		.d(n3378), .sdi(n1930), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__29__slave ( .q(_RegFile_11__29), .qb(n1931),
		.d(_RegFile_reg_11__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__2__master ( .q(_RegFile_reg_11__2__m2s), .qb(),
		.d(n3351), .sdi(n4279), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__2__slave ( .q(_RegFile_11__2), .qb(n4278), .d(_RegFile_reg_11__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__30__master ( .q(_RegFile_reg_11__30__m2s), .qb(),
		.d(n3379), .sdi(n1931), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__30__slave ( .q(_RegFile_11__30), .qb(n1932),
		.d(_RegFile_reg_11__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__31__master ( .q(_RegFile_reg_11__31__m2s), .qb(),
		.d(n3380), .sdi(n1932), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__31__slave ( .q(_RegFile_11__31), .qb(n1933),
		.d(_RegFile_reg_11__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__3__master ( .q(_RegFile_reg_11__3__m2s), .qb(),
		.d(n3352), .sdi(n4278), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__3__slave ( .q(_RegFile_11__3), .qb(n4277), .d(_RegFile_reg_11__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__4__master ( .q(_RegFile_reg_11__4__m2s), .qb(),
		.d(n3353), .sdi(n4277), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__4__slave ( .q(_RegFile_11__4), .qb(n4276), .d(_RegFile_reg_11__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__5__master ( .q(_RegFile_reg_11__5__m2s), .qb(),
		.d(n3354), .sdi(n4276), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__5__slave ( .q(_RegFile_11__5), .qb(n4275), .d(_RegFile_reg_11__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__6__master ( .q(_RegFile_reg_11__6__m2s), .qb(),
		.d(n3355), .sdi(n4275), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__6__slave ( .q(_RegFile_11__6), .qb(n4274), .d(_RegFile_reg_11__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__7__master ( .q(_RegFile_reg_11__7__m2s), .qb(),
		.d(n3356), .sdi(n4274), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__7__slave ( .q(_RegFile_11__7), .qb(n4273), .d(_RegFile_reg_11__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__8__master ( .q(_RegFile_reg_11__8__m2s), .qb(),
		.d(n3357), .sdi(n4273), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__8__slave ( .q(_RegFile_11__8), .qb(n1934), .d(_RegFile_reg_11__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_11__9__master ( .q(_RegFile_reg_11__9__m2s), .qb(),
		.d(n3358), .sdi(n1934), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_11__9__slave ( .q(_RegFile_11__9), .qb(n1935), .d(_RegFile_reg_11__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__0__master ( .q(_RegFile_reg_12__0__m2s), .qb(),
		.d(n3317), .sdi(n1933), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n958),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__0__slave ( .q(_RegFile_12__0), .qb(n4272), .d(_RegFile_reg_12__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n958), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__10__master ( .q(_RegFile_reg_12__10__m2s), .qb(),
		.d(n3327), .sdi(n1959), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__10__slave ( .q(_RegFile_12__10), .qb(n1936),
		.d(_RegFile_reg_12__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__11__master ( .q(_RegFile_reg_12__11__m2s), .qb(),
		.d(n3328), .sdi(n1936), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__11__slave ( .q(_RegFile_12__11), .qb(n1937),
		.d(_RegFile_reg_12__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__12__master ( .q(_RegFile_reg_12__12__m2s), .qb(),
		.d(n3329), .sdi(n1937), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__12__slave ( .q(_RegFile_12__12), .qb(n1938),
		.d(_RegFile_reg_12__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__13__master ( .q(_RegFile_reg_12__13__m2s), .qb(),
		.d(n3330), .sdi(n1938), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__13__slave ( .q(_RegFile_12__13), .qb(n1939),
		.d(_RegFile_reg_12__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__14__master ( .q(_RegFile_reg_12__14__m2s), .qb(),
		.d(n3331), .sdi(n1939), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__14__slave ( .q(_RegFile_12__14), .qb(n1940),
		.d(_RegFile_reg_12__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__15__master ( .q(_RegFile_reg_12__15__m2s), .qb(),
		.d(n3332), .sdi(n1940), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__15__slave ( .q(_RegFile_12__15), .qb(n1941),
		.d(_RegFile_reg_12__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__16__master ( .q(_RegFile_reg_12__16__m2s), .qb(),
		.d(n3333), .sdi(n1941), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__16__slave ( .q(_RegFile_12__16), .qb(n1942),
		.d(_RegFile_reg_12__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__17__master ( .q(_RegFile_reg_12__17__m2s), .qb(),
		.d(n3334), .sdi(n1942), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__17__slave ( .q(_RegFile_12__17), .qb(n1943),
		.d(_RegFile_reg_12__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__18__master ( .q(_RegFile_reg_12__18__m2s), .qb(),
		.d(n3335), .sdi(n1943), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__18__slave ( .q(_RegFile_12__18), .qb(n1944),
		.d(_RegFile_reg_12__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__19__master ( .q(_RegFile_reg_12__19__m2s), .qb(),
		.d(n3336), .sdi(n1944), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__19__slave ( .q(_RegFile_12__19), .qb(n1945),
		.d(_RegFile_reg_12__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__1__master ( .q(_RegFile_reg_12__1__m2s), .qb(),
		.d(n3318), .sdi(n4272), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__1__slave ( .q(_RegFile_12__1), .qb(n4271), .d(_RegFile_reg_12__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__20__master ( .q(_RegFile_reg_12__20__m2s), .qb(),
		.d(n3337), .sdi(n1945), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__20__slave ( .q(_RegFile_12__20), .qb(n1946),
		.d(_RegFile_reg_12__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__21__master ( .q(_RegFile_reg_12__21__m2s), .qb(),
		.d(n3338), .sdi(n1946), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__21__slave ( .q(_RegFile_12__21), .qb(n1947),
		.d(_RegFile_reg_12__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__22__master ( .q(_RegFile_reg_12__22__m2s), .qb(),
		.d(n3339), .sdi(n1947), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__22__slave ( .q(_RegFile_12__22), .qb(n1948),
		.d(_RegFile_reg_12__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__23__master ( .q(_RegFile_reg_12__23__m2s), .qb(),
		.d(n3340), .sdi(n1948), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__23__slave ( .q(_RegFile_12__23), .qb(n1949),
		.d(_RegFile_reg_12__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__24__master ( .q(_RegFile_reg_12__24__m2s), .qb(),
		.d(n3341), .sdi(n1949), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__24__slave ( .q(_RegFile_12__24), .qb(n1950),
		.d(_RegFile_reg_12__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__25__master ( .q(_RegFile_reg_12__25__m2s), .qb(),
		.d(n3342), .sdi(n1950), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__25__slave ( .q(_RegFile_12__25), .qb(n1951),
		.d(_RegFile_reg_12__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__26__master ( .q(_RegFile_reg_12__26__m2s), .qb(),
		.d(n3343), .sdi(n1951), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__26__slave ( .q(_RegFile_12__26), .qb(n1952),
		.d(_RegFile_reg_12__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__27__master ( .q(_RegFile_reg_12__27__m2s), .qb(),
		.d(n3344), .sdi(n1952), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__27__slave ( .q(_RegFile_12__27), .qb(n1953),
		.d(_RegFile_reg_12__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__28__master ( .q(_RegFile_reg_12__28__m2s), .qb(),
		.d(n3345), .sdi(n1953), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__28__slave ( .q(_RegFile_12__28), .qb(n1954),
		.d(_RegFile_reg_12__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__29__master ( .q(_RegFile_reg_12__29__m2s), .qb(),
		.d(n3346), .sdi(n1954), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__29__slave ( .q(_RegFile_12__29), .qb(n1955),
		.d(_RegFile_reg_12__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__2__master ( .q(_RegFile_reg_12__2__m2s), .qb(),
		.d(n3319), .sdi(n4271), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__2__slave ( .q(_RegFile_12__2), .qb(n4270), .d(_RegFile_reg_12__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__30__master ( .q(_RegFile_reg_12__30__m2s), .qb(),
		.d(n3347), .sdi(n1955), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__30__slave ( .q(_RegFile_12__30), .qb(n1956),
		.d(_RegFile_reg_12__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__31__master ( .q(_RegFile_reg_12__31__m2s), .qb(),
		.d(n3348), .sdi(n1956), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__31__slave ( .q(_RegFile_12__31), .qb(n1957),
		.d(_RegFile_reg_12__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__3__master ( .q(_RegFile_reg_12__3__m2s), .qb(),
		.d(n3320), .sdi(n4270), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__3__slave ( .q(_RegFile_12__3), .qb(n4269), .d(_RegFile_reg_12__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__4__master ( .q(_RegFile_reg_12__4__m2s), .qb(),
		.d(n3321), .sdi(n4269), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__4__slave ( .q(_RegFile_12__4), .qb(n4268), .d(_RegFile_reg_12__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__5__master ( .q(_RegFile_reg_12__5__m2s), .qb(),
		.d(n3322), .sdi(n4268), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__5__slave ( .q(_RegFile_12__5), .qb(n4267), .d(_RegFile_reg_12__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__6__master ( .q(_RegFile_reg_12__6__m2s), .qb(),
		.d(n3323), .sdi(n4267), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__6__slave ( .q(_RegFile_12__6), .qb(n4266), .d(_RegFile_reg_12__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__7__master ( .q(_RegFile_reg_12__7__m2s), .qb(),
		.d(n3324), .sdi(n4266), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__7__slave ( .q(_RegFile_12__7), .qb(n4265), .d(_RegFile_reg_12__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__8__master ( .q(_RegFile_reg_12__8__m2s), .qb(),
		.d(n3325), .sdi(n4265), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n959),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__8__slave ( .q(_RegFile_12__8), .qb(n1958), .d(_RegFile_reg_12__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n959), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_12__9__master ( .q(_RegFile_reg_12__9__m2s), .qb(),
		.d(n3326), .sdi(n1958), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_12__9__slave ( .q(_RegFile_12__9), .qb(n1959), .d(_RegFile_reg_12__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__0__master ( .q(_RegFile_reg_13__0__m2s), .qb(),
		.d(n3285), .sdi(n1957), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__0__slave ( .q(_RegFile_13__0), .qb(n4264), .d(_RegFile_reg_13__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__10__master ( .q(_RegFile_reg_13__10__m2s), .qb(),
		.d(n3295), .sdi(n1983), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__10__slave ( .q(_RegFile_13__10), .qb(n1960),
		.d(_RegFile_reg_13__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__11__master ( .q(_RegFile_reg_13__11__m2s), .qb(),
		.d(n3296), .sdi(n1960), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__11__slave ( .q(_RegFile_13__11), .qb(n1961),
		.d(_RegFile_reg_13__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__12__master ( .q(_RegFile_reg_13__12__m2s), .qb(),
		.d(n3297), .sdi(n1961), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__12__slave ( .q(_RegFile_13__12), .qb(n1962),
		.d(_RegFile_reg_13__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__13__master ( .q(_RegFile_reg_13__13__m2s), .qb(),
		.d(n3298), .sdi(n1962), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__13__slave ( .q(_RegFile_13__13), .qb(n1963),
		.d(_RegFile_reg_13__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__14__master ( .q(_RegFile_reg_13__14__m2s), .qb(),
		.d(n3299), .sdi(n1963), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__14__slave ( .q(_RegFile_13__14), .qb(n1964),
		.d(_RegFile_reg_13__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__15__master ( .q(_RegFile_reg_13__15__m2s), .qb(),
		.d(n3300), .sdi(n1964), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__15__slave ( .q(_RegFile_13__15), .qb(n1965),
		.d(_RegFile_reg_13__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__16__master ( .q(_RegFile_reg_13__16__m2s), .qb(),
		.d(n3301), .sdi(n1965), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__16__slave ( .q(_RegFile_13__16), .qb(n1966),
		.d(_RegFile_reg_13__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__17__master ( .q(_RegFile_reg_13__17__m2s), .qb(),
		.d(n3302), .sdi(n1966), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__17__slave ( .q(_RegFile_13__17), .qb(n1967),
		.d(_RegFile_reg_13__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__18__master ( .q(_RegFile_reg_13__18__m2s), .qb(),
		.d(n3303), .sdi(n1967), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__18__slave ( .q(_RegFile_13__18), .qb(n1968),
		.d(_RegFile_reg_13__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__19__master ( .q(_RegFile_reg_13__19__m2s), .qb(),
		.d(n3304), .sdi(n1968), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__19__slave ( .q(_RegFile_13__19), .qb(n1969),
		.d(_RegFile_reg_13__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__1__master ( .q(_RegFile_reg_13__1__m2s), .qb(),
		.d(n3286), .sdi(n4264), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__1__slave ( .q(_RegFile_13__1), .qb(n4263), .d(_RegFile_reg_13__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__20__master ( .q(_RegFile_reg_13__20__m2s), .qb(),
		.d(n3305), .sdi(n1969), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n946),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__20__slave ( .q(_RegFile_13__20), .qb(n1970),
		.d(_RegFile_reg_13__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n946), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__21__master ( .q(_RegFile_reg_13__21__m2s), .qb(),
		.d(n3306), .sdi(n1970), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__21__slave ( .q(_RegFile_13__21), .qb(n1971),
		.d(_RegFile_reg_13__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__22__master ( .q(_RegFile_reg_13__22__m2s), .qb(),
		.d(n3307), .sdi(n1971), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__22__slave ( .q(_RegFile_13__22), .qb(n1972),
		.d(_RegFile_reg_13__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__23__master ( .q(_RegFile_reg_13__23__m2s), .qb(),
		.d(n3308), .sdi(n1972), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__23__slave ( .q(_RegFile_13__23), .qb(n1973),
		.d(_RegFile_reg_13__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__24__master ( .q(_RegFile_reg_13__24__m2s), .qb(),
		.d(n3309), .sdi(n1973), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__24__slave ( .q(_RegFile_13__24), .qb(n1974),
		.d(_RegFile_reg_13__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__25__master ( .q(_RegFile_reg_13__25__m2s), .qb(),
		.d(n3310), .sdi(n1974), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__25__slave ( .q(_RegFile_13__25), .qb(n1975),
		.d(_RegFile_reg_13__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__26__master ( .q(_RegFile_reg_13__26__m2s), .qb(),
		.d(n3311), .sdi(n1975), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__26__slave ( .q(_RegFile_13__26), .qb(n1976),
		.d(_RegFile_reg_13__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__27__master ( .q(_RegFile_reg_13__27__m2s), .qb(),
		.d(n3312), .sdi(n1976), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__27__slave ( .q(_RegFile_13__27), .qb(n1977),
		.d(_RegFile_reg_13__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__28__master ( .q(_RegFile_reg_13__28__m2s), .qb(),
		.d(n3313), .sdi(n1977), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__28__slave ( .q(_RegFile_13__28), .qb(n1978),
		.d(_RegFile_reg_13__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__29__master ( .q(_RegFile_reg_13__29__m2s), .qb(),
		.d(n3314), .sdi(n1978), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__29__slave ( .q(_RegFile_13__29), .qb(n1979),
		.d(_RegFile_reg_13__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__2__master ( .q(_RegFile_reg_13__2__m2s), .qb(),
		.d(n3287), .sdi(n4263), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__2__slave ( .q(_RegFile_13__2), .qb(n4262), .d(_RegFile_reg_13__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__30__master ( .q(_RegFile_reg_13__30__m2s), .qb(),
		.d(n3315), .sdi(n1979), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__30__slave ( .q(_RegFile_13__30), .qb(n1980),
		.d(_RegFile_reg_13__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__31__master ( .q(_RegFile_reg_13__31__m2s), .qb(),
		.d(n3316), .sdi(n1980), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__31__slave ( .q(_RegFile_13__31), .qb(n1981),
		.d(_RegFile_reg_13__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__3__master ( .q(_RegFile_reg_13__3__m2s), .qb(),
		.d(n3288), .sdi(n4262), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__3__slave ( .q(_RegFile_13__3), .qb(n4261), .d(_RegFile_reg_13__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__4__master ( .q(_RegFile_reg_13__4__m2s), .qb(),
		.d(n3289), .sdi(n4261), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__4__slave ( .q(_RegFile_13__4), .qb(n4260), .d(_RegFile_reg_13__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__5__master ( .q(_RegFile_reg_13__5__m2s), .qb(),
		.d(n3290), .sdi(n4260), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__5__slave ( .q(_RegFile_13__5), .qb(n4259), .d(_RegFile_reg_13__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__6__master ( .q(_RegFile_reg_13__6__m2s), .qb(),
		.d(n3291), .sdi(n4259), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__6__slave ( .q(_RegFile_13__6), .qb(n4258), .d(_RegFile_reg_13__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__7__master ( .q(_RegFile_reg_13__7__m2s), .qb(),
		.d(n3292), .sdi(n4258), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__7__slave ( .q(_RegFile_13__7), .qb(n4257), .d(_RegFile_reg_13__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__8__master ( .q(_RegFile_reg_13__8__m2s), .qb(),
		.d(n3293), .sdi(n4257), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__8__slave ( .q(_RegFile_13__8), .qb(n1982), .d(_RegFile_reg_13__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_13__9__master ( .q(_RegFile_reg_13__9__m2s), .qb(),
		.d(n3294), .sdi(n1982), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_13__9__slave ( .q(_RegFile_13__9), .qb(n1983), .d(_RegFile_reg_13__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__0__master ( .q(_RegFile_reg_14__0__m2s), .qb(),
		.d(n3253), .sdi(n1981), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__0__slave ( .q(_RegFile_14__0), .qb(n4256), .d(_RegFile_reg_14__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__10__master ( .q(_RegFile_reg_14__10__m2s), .qb(),
		.d(n3263), .sdi(n2007), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__10__slave ( .q(_RegFile_14__10), .qb(n1984),
		.d(_RegFile_reg_14__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__11__master ( .q(_RegFile_reg_14__11__m2s), .qb(),
		.d(n3264), .sdi(n1984), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__11__slave ( .q(_RegFile_14__11), .qb(n1985),
		.d(_RegFile_reg_14__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__12__master ( .q(_RegFile_reg_14__12__m2s), .qb(),
		.d(n3265), .sdi(n1985), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__12__slave ( .q(_RegFile_14__12), .qb(n1986),
		.d(_RegFile_reg_14__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__13__master ( .q(_RegFile_reg_14__13__m2s), .qb(),
		.d(n3266), .sdi(n1986), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__13__slave ( .q(_RegFile_14__13), .qb(n1987),
		.d(_RegFile_reg_14__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__14__master ( .q(_RegFile_reg_14__14__m2s), .qb(),
		.d(n3267), .sdi(n1987), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__14__slave ( .q(_RegFile_14__14), .qb(n1988),
		.d(_RegFile_reg_14__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__15__master ( .q(_RegFile_reg_14__15__m2s), .qb(),
		.d(n3268), .sdi(n1988), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__15__slave ( .q(_RegFile_14__15), .qb(n1989),
		.d(_RegFile_reg_14__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__16__master ( .q(_RegFile_reg_14__16__m2s), .qb(),
		.d(n3269), .sdi(n1989), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__16__slave ( .q(_RegFile_14__16), .qb(n1990),
		.d(_RegFile_reg_14__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__17__master ( .q(_RegFile_reg_14__17__m2s), .qb(),
		.d(n3270), .sdi(n1990), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__17__slave ( .q(_RegFile_14__17), .qb(n1991),
		.d(_RegFile_reg_14__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__18__master ( .q(_RegFile_reg_14__18__m2s), .qb(),
		.d(n3271), .sdi(n1991), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__18__slave ( .q(_RegFile_14__18), .qb(n1992),
		.d(_RegFile_reg_14__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__19__master ( .q(_RegFile_reg_14__19__m2s), .qb(),
		.d(n3272), .sdi(n1992), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__19__slave ( .q(_RegFile_14__19), .qb(n1993),
		.d(_RegFile_reg_14__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__1__master ( .q(_RegFile_reg_14__1__m2s), .qb(),
		.d(n3254), .sdi(n4256), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n945),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__1__slave ( .q(_RegFile_14__1), .qb(n4255), .d(_RegFile_reg_14__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n945), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__20__master ( .q(_RegFile_reg_14__20__m2s), .qb(),
		.d(n3273), .sdi(n1993), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__20__slave ( .q(_RegFile_14__20), .qb(n1994),
		.d(_RegFile_reg_14__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__21__master ( .q(_RegFile_reg_14__21__m2s), .qb(),
		.d(n3274), .sdi(n1994), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__21__slave ( .q(_RegFile_14__21), .qb(n1995),
		.d(_RegFile_reg_14__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__22__master ( .q(_RegFile_reg_14__22__m2s), .qb(),
		.d(n3275), .sdi(n1995), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__22__slave ( .q(_RegFile_14__22), .qb(n1996),
		.d(_RegFile_reg_14__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__23__master ( .q(_RegFile_reg_14__23__m2s), .qb(),
		.d(n3276), .sdi(n1996), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__23__slave ( .q(_RegFile_14__23), .qb(n1997),
		.d(_RegFile_reg_14__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__24__master ( .q(_RegFile_reg_14__24__m2s), .qb(),
		.d(n3277), .sdi(n1997), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__24__slave ( .q(_RegFile_14__24), .qb(n1998),
		.d(_RegFile_reg_14__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__25__master ( .q(_RegFile_reg_14__25__m2s), .qb(),
		.d(n3278), .sdi(n1998), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__25__slave ( .q(_RegFile_14__25), .qb(n1999),
		.d(_RegFile_reg_14__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__26__master ( .q(_RegFile_reg_14__26__m2s), .qb(),
		.d(n3279), .sdi(n1999), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__26__slave ( .q(_RegFile_14__26), .qb(n2000),
		.d(_RegFile_reg_14__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__27__master ( .q(_RegFile_reg_14__27__m2s), .qb(),
		.d(n3280), .sdi(n2000), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__27__slave ( .q(_RegFile_14__27), .qb(n2001),
		.d(_RegFile_reg_14__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__28__master ( .q(_RegFile_reg_14__28__m2s), .qb(),
		.d(n3281), .sdi(n2001), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__28__slave ( .q(_RegFile_14__28), .qb(n2002),
		.d(_RegFile_reg_14__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__29__master ( .q(_RegFile_reg_14__29__m2s), .qb(),
		.d(n3282), .sdi(n2002), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__29__slave ( .q(_RegFile_14__29), .qb(n2003),
		.d(_RegFile_reg_14__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__2__master ( .q(_RegFile_reg_14__2__m2s), .qb(),
		.d(n3255), .sdi(n4255), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__2__slave ( .q(_RegFile_14__2), .qb(n4254), .d(_RegFile_reg_14__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__30__master ( .q(_RegFile_reg_14__30__m2s), .qb(),
		.d(n3283), .sdi(n2003), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__30__slave ( .q(_RegFile_14__30), .qb(n2004),
		.d(_RegFile_reg_14__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__31__master ( .q(_RegFile_reg_14__31__m2s), .qb(),
		.d(n3284), .sdi(n2004), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__31__slave ( .q(_RegFile_14__31), .qb(n2005),
		.d(_RegFile_reg_14__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__3__master ( .q(_RegFile_reg_14__3__m2s), .qb(),
		.d(n3256), .sdi(n4254), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__3__slave ( .q(_RegFile_14__3), .qb(n4253), .d(_RegFile_reg_14__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__4__master ( .q(_RegFile_reg_14__4__m2s), .qb(),
		.d(n3257), .sdi(n4253), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__4__slave ( .q(_RegFile_14__4), .qb(n4252), .d(_RegFile_reg_14__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__5__master ( .q(_RegFile_reg_14__5__m2s), .qb(),
		.d(n3258), .sdi(n4252), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__5__slave ( .q(_RegFile_14__5), .qb(n4251), .d(_RegFile_reg_14__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__6__master ( .q(_RegFile_reg_14__6__m2s), .qb(),
		.d(n3259), .sdi(n4251), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__6__slave ( .q(_RegFile_14__6), .qb(n4250), .d(_RegFile_reg_14__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__7__master ( .q(_RegFile_reg_14__7__m2s), .qb(),
		.d(n3260), .sdi(n4250), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__7__slave ( .q(_RegFile_14__7), .qb(n4249), .d(_RegFile_reg_14__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__8__master ( .q(_RegFile_reg_14__8__m2s), .qb(),
		.d(n3261), .sdi(n4249), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__8__slave ( .q(_RegFile_14__8), .qb(n2006), .d(_RegFile_reg_14__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_14__9__master ( .q(_RegFile_reg_14__9__m2s), .qb(),
		.d(n3262), .sdi(n2006), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_14__9__slave ( .q(_RegFile_14__9), .qb(n2007), .d(_RegFile_reg_14__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__0__master ( .q(_RegFile_reg_15__0__m2s), .qb(),
		.d(n3221), .sdi(n2005), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__0__slave ( .q(_RegFile_15__0), .qb(n4248), .d(_RegFile_reg_15__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__10__master ( .q(_RegFile_reg_15__10__m2s), .qb(),
		.d(n3231), .sdi(n2031), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__10__slave ( .q(_RegFile_15__10), .qb(n2008),
		.d(_RegFile_reg_15__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__11__master ( .q(_RegFile_reg_15__11__m2s), .qb(),
		.d(n3232), .sdi(n2008), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__11__slave ( .q(_RegFile_15__11), .qb(n2009),
		.d(_RegFile_reg_15__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__12__master ( .q(_RegFile_reg_15__12__m2s), .qb(),
		.d(n3233), .sdi(n2009), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__12__slave ( .q(_RegFile_15__12), .qb(n2010),
		.d(_RegFile_reg_15__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__13__master ( .q(_RegFile_reg_15__13__m2s), .qb(),
		.d(n3234), .sdi(n2010), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__13__slave ( .q(_RegFile_15__13), .qb(n2011),
		.d(_RegFile_reg_15__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__14__master ( .q(_RegFile_reg_15__14__m2s), .qb(),
		.d(n3235), .sdi(n2011), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__14__slave ( .q(_RegFile_15__14), .qb(n2012),
		.d(_RegFile_reg_15__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__15__master ( .q(_RegFile_reg_15__15__m2s), .qb(),
		.d(n3236), .sdi(n2012), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__15__slave ( .q(_RegFile_15__15), .qb(n2013),
		.d(_RegFile_reg_15__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__16__master ( .q(_RegFile_reg_15__16__m2s), .qb(),
		.d(n3237), .sdi(n2013), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__16__slave ( .q(_RegFile_15__16), .qb(n2014),
		.d(_RegFile_reg_15__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__17__master ( .q(_RegFile_reg_15__17__m2s), .qb(),
		.d(n3238), .sdi(n2014), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__17__slave ( .q(_RegFile_15__17), .qb(n2015),
		.d(_RegFile_reg_15__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__18__master ( .q(_RegFile_reg_15__18__m2s), .qb(),
		.d(n3239), .sdi(n2015), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__18__slave ( .q(_RegFile_15__18), .qb(n2016),
		.d(_RegFile_reg_15__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__19__master ( .q(_RegFile_reg_15__19__m2s), .qb(),
		.d(n3240), .sdi(n2016), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__19__slave ( .q(_RegFile_15__19), .qb(n2017),
		.d(_RegFile_reg_15__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__1__master ( .q(_RegFile_reg_15__1__m2s), .qb(),
		.d(n3222), .sdi(n4248), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__1__slave ( .q(_RegFile_15__1), .qb(n4247), .d(_RegFile_reg_15__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__20__master ( .q(_RegFile_reg_15__20__m2s), .qb(),
		.d(n3241), .sdi(n2017), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__20__slave ( .q(_RegFile_15__20), .qb(n2018),
		.d(_RegFile_reg_15__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__21__master ( .q(_RegFile_reg_15__21__m2s), .qb(),
		.d(n3242), .sdi(n2018), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__21__slave ( .q(_RegFile_15__21), .qb(n2019),
		.d(_RegFile_reg_15__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__22__master ( .q(_RegFile_reg_15__22__m2s), .qb(),
		.d(n3243), .sdi(n2019), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__22__slave ( .q(_RegFile_15__22), .qb(n2020),
		.d(_RegFile_reg_15__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__23__master ( .q(_RegFile_reg_15__23__m2s), .qb(),
		.d(n3244), .sdi(n2020), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__23__slave ( .q(_RegFile_15__23), .qb(n2021),
		.d(_RegFile_reg_15__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__24__master ( .q(_RegFile_reg_15__24__m2s), .qb(),
		.d(n3245), .sdi(n2021), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__24__slave ( .q(_RegFile_15__24), .qb(n2022),
		.d(_RegFile_reg_15__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__25__master ( .q(_RegFile_reg_15__25__m2s), .qb(),
		.d(n3246), .sdi(n2022), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__25__slave ( .q(_RegFile_15__25), .qb(n2023),
		.d(_RegFile_reg_15__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__26__master ( .q(_RegFile_reg_15__26__m2s), .qb(),
		.d(n3247), .sdi(n2023), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__26__slave ( .q(_RegFile_15__26), .qb(n2024),
		.d(_RegFile_reg_15__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__27__master ( .q(_RegFile_reg_15__27__m2s), .qb(),
		.d(n3248), .sdi(n2024), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__27__slave ( .q(_RegFile_15__27), .qb(n2025),
		.d(_RegFile_reg_15__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__28__master ( .q(_RegFile_reg_15__28__m2s), .qb(),
		.d(n3249), .sdi(n2025), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__28__slave ( .q(_RegFile_15__28), .qb(n2026),
		.d(_RegFile_reg_15__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__29__master ( .q(_RegFile_reg_15__29__m2s), .qb(),
		.d(n3250), .sdi(n2026), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__29__slave ( .q(_RegFile_15__29), .qb(n2027),
		.d(_RegFile_reg_15__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__2__master ( .q(_RegFile_reg_15__2__m2s), .qb(),
		.d(n3223), .sdi(n4247), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__2__slave ( .q(_RegFile_15__2), .qb(n4246), .d(_RegFile_reg_15__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__30__master ( .q(_RegFile_reg_15__30__m2s), .qb(),
		.d(n3251), .sdi(n2027), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__30__slave ( .q(_RegFile_15__30), .qb(n2028),
		.d(_RegFile_reg_15__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__31__master ( .q(_RegFile_reg_15__31__m2s), .qb(),
		.d(n3252), .sdi(n2028), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__31__slave ( .q(_RegFile_15__31), .qb(n2029),
		.d(_RegFile_reg_15__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__3__master ( .q(_RegFile_reg_15__3__m2s), .qb(),
		.d(n3224), .sdi(n4246), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__3__slave ( .q(_RegFile_15__3), .qb(n4245), .d(_RegFile_reg_15__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__4__master ( .q(_RegFile_reg_15__4__m2s), .qb(),
		.d(n3225), .sdi(n4245), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__4__slave ( .q(_RegFile_15__4), .qb(n4244), .d(_RegFile_reg_15__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__5__master ( .q(_RegFile_reg_15__5__m2s), .qb(),
		.d(n3226), .sdi(n4244), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__5__slave ( .q(_RegFile_15__5), .qb(n4243), .d(_RegFile_reg_15__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__6__master ( .q(_RegFile_reg_15__6__m2s), .qb(),
		.d(n3227), .sdi(n4243), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__6__slave ( .q(_RegFile_15__6), .qb(n4242), .d(_RegFile_reg_15__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__7__master ( .q(_RegFile_reg_15__7__m2s), .qb(),
		.d(n3228), .sdi(n4242), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__7__slave ( .q(_RegFile_15__7), .qb(n4241), .d(_RegFile_reg_15__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__8__master ( .q(_RegFile_reg_15__8__m2s), .qb(),
		.d(n3229), .sdi(n4241), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__8__slave ( .q(_RegFile_15__8), .qb(n2030), .d(_RegFile_reg_15__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_15__9__master ( .q(_RegFile_reg_15__9__m2s), .qb(),
		.d(n3230), .sdi(n2030), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_15__9__slave ( .q(_RegFile_15__9), .qb(n2031), .d(_RegFile_reg_15__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__0__master ( .q(_RegFile_reg_16__0__m2s), .qb(),
		.d(n3189), .sdi(n2029), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__0__slave ( .q(_RegFile_16__0), .qb(n4240), .d(_RegFile_reg_16__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__10__master ( .q(_RegFile_reg_16__10__m2s), .qb(),
		.d(n3199), .sdi(n2055), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__10__slave ( .q(_RegFile_16__10), .qb(n2032),
		.d(_RegFile_reg_16__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__11__master ( .q(_RegFile_reg_16__11__m2s), .qb(),
		.d(n3200), .sdi(n2032), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__11__slave ( .q(_RegFile_16__11), .qb(n2033),
		.d(_RegFile_reg_16__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__12__master ( .q(_RegFile_reg_16__12__m2s), .qb(),
		.d(n3201), .sdi(n2033), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__12__slave ( .q(_RegFile_16__12), .qb(n2034),
		.d(_RegFile_reg_16__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__13__master ( .q(_RegFile_reg_16__13__m2s), .qb(),
		.d(n3202), .sdi(n2034), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__13__slave ( .q(_RegFile_16__13), .qb(n2035),
		.d(_RegFile_reg_16__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__14__master ( .q(_RegFile_reg_16__14__m2s), .qb(),
		.d(n3203), .sdi(n2035), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__14__slave ( .q(_RegFile_16__14), .qb(n2036),
		.d(_RegFile_reg_16__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__15__master ( .q(_RegFile_reg_16__15__m2s), .qb(),
		.d(n3204), .sdi(n2036), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__15__slave ( .q(_RegFile_16__15), .qb(n2037),
		.d(_RegFile_reg_16__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__16__master ( .q(_RegFile_reg_16__16__m2s), .qb(),
		.d(n3205), .sdi(n2037), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__16__slave ( .q(_RegFile_16__16), .qb(n2038),
		.d(_RegFile_reg_16__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__17__master ( .q(_RegFile_reg_16__17__m2s), .qb(),
		.d(n3206), .sdi(n2038), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__17__slave ( .q(_RegFile_16__17), .qb(n2039),
		.d(_RegFile_reg_16__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__18__master ( .q(_RegFile_reg_16__18__m2s), .qb(),
		.d(n3207), .sdi(n2039), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__18__slave ( .q(_RegFile_16__18), .qb(n2040),
		.d(_RegFile_reg_16__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__19__master ( .q(_RegFile_reg_16__19__m2s), .qb(),
		.d(n3208), .sdi(n2040), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__19__slave ( .q(_RegFile_16__19), .qb(n2041),
		.d(_RegFile_reg_16__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__1__master ( .q(_RegFile_reg_16__1__m2s), .qb(),
		.d(n3190), .sdi(n4240), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n944),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__1__slave ( .q(_RegFile_16__1), .qb(n4239), .d(_RegFile_reg_16__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n944), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__20__master ( .q(_RegFile_reg_16__20__m2s), .qb(),
		.d(n3209), .sdi(n2041), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__20__slave ( .q(_RegFile_16__20), .qb(n2042),
		.d(_RegFile_reg_16__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__21__master ( .q(_RegFile_reg_16__21__m2s), .qb(),
		.d(n3210), .sdi(n2042), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__21__slave ( .q(_RegFile_16__21), .qb(n2043),
		.d(_RegFile_reg_16__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__22__master ( .q(_RegFile_reg_16__22__m2s), .qb(),
		.d(n3211), .sdi(n2043), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__22__slave ( .q(_RegFile_16__22), .qb(n2044),
		.d(_RegFile_reg_16__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__23__master ( .q(_RegFile_reg_16__23__m2s), .qb(),
		.d(n3212), .sdi(n2044), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__23__slave ( .q(_RegFile_16__23), .qb(n2045),
		.d(_RegFile_reg_16__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__24__master ( .q(_RegFile_reg_16__24__m2s), .qb(),
		.d(n3213), .sdi(n2045), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__24__slave ( .q(_RegFile_16__24), .qb(n2046),
		.d(_RegFile_reg_16__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__25__master ( .q(_RegFile_reg_16__25__m2s), .qb(),
		.d(n3214), .sdi(n2046), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__25__slave ( .q(_RegFile_16__25), .qb(n2047),
		.d(_RegFile_reg_16__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__26__master ( .q(_RegFile_reg_16__26__m2s), .qb(),
		.d(n3215), .sdi(n2047), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__26__slave ( .q(_RegFile_16__26), .qb(n2048),
		.d(_RegFile_reg_16__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__27__master ( .q(_RegFile_reg_16__27__m2s), .qb(),
		.d(n3216), .sdi(n2048), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__27__slave ( .q(_RegFile_16__27), .qb(n2049),
		.d(_RegFile_reg_16__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__28__master ( .q(_RegFile_reg_16__28__m2s), .qb(),
		.d(n3217), .sdi(n2049), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__28__slave ( .q(_RegFile_16__28), .qb(n2050),
		.d(_RegFile_reg_16__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__29__master ( .q(_RegFile_reg_16__29__m2s), .qb(),
		.d(n3218), .sdi(n2050), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__29__slave ( .q(_RegFile_16__29), .qb(n2051),
		.d(_RegFile_reg_16__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__2__master ( .q(_RegFile_reg_16__2__m2s), .qb(),
		.d(n3191), .sdi(n4239), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n960),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__2__slave ( .q(_RegFile_16__2), .qb(n4238), .d(_RegFile_reg_16__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n960), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__30__master ( .q(_RegFile_reg_16__30__m2s), .qb(),
		.d(n3219), .sdi(n2051), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__30__slave ( .q(_RegFile_16__30), .qb(n2052),
		.d(_RegFile_reg_16__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__31__master ( .q(_RegFile_reg_16__31__m2s), .qb(),
		.d(n3220), .sdi(n2052), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__31__slave ( .q(_RegFile_16__31), .qb(n2053),
		.d(_RegFile_reg_16__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__3__master ( .q(_RegFile_reg_16__3__m2s), .qb(),
		.d(n3192), .sdi(n4238), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__3__slave ( .q(_RegFile_16__3), .qb(n4237), .d(_RegFile_reg_16__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__4__master ( .q(_RegFile_reg_16__4__m2s), .qb(),
		.d(n3193), .sdi(n4237), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__4__slave ( .q(_RegFile_16__4), .qb(n4236), .d(_RegFile_reg_16__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__5__master ( .q(_RegFile_reg_16__5__m2s), .qb(),
		.d(n3194), .sdi(n4236), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__5__slave ( .q(_RegFile_16__5), .qb(n4235), .d(_RegFile_reg_16__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__6__master ( .q(_RegFile_reg_16__6__m2s), .qb(),
		.d(n3195), .sdi(n4235), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__6__slave ( .q(_RegFile_16__6), .qb(n4234), .d(_RegFile_reg_16__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__7__master ( .q(_RegFile_reg_16__7__m2s), .qb(),
		.d(n3196), .sdi(n4234), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__7__slave ( .q(_RegFile_16__7), .qb(n4233), .d(_RegFile_reg_16__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__8__master ( .q(_RegFile_reg_16__8__m2s), .qb(),
		.d(n3197), .sdi(n4233), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__8__slave ( .q(_RegFile_16__8), .qb(n2054), .d(_RegFile_reg_16__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_16__9__master ( .q(_RegFile_reg_16__9__m2s), .qb(),
		.d(n3198), .sdi(n2054), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_16__9__slave ( .q(_RegFile_16__9), .qb(n2055), .d(_RegFile_reg_16__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__0__master ( .q(_RegFile_reg_17__0__m2s), .qb(),
		.d(n3157), .sdi(n2053), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__0__slave ( .q(_RegFile_17__0), .qb(n4232), .d(_RegFile_reg_17__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__10__master ( .q(_RegFile_reg_17__10__m2s), .qb(),
		.d(n3167), .sdi(n2079), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__10__slave ( .q(_RegFile_17__10), .qb(n2056),
		.d(_RegFile_reg_17__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__11__master ( .q(_RegFile_reg_17__11__m2s), .qb(),
		.d(n3168), .sdi(n2056), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__11__slave ( .q(_RegFile_17__11), .qb(n2057),
		.d(_RegFile_reg_17__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__12__master ( .q(_RegFile_reg_17__12__m2s), .qb(),
		.d(n3169), .sdi(n2057), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__12__slave ( .q(_RegFile_17__12), .qb(n2058),
		.d(_RegFile_reg_17__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__13__master ( .q(_RegFile_reg_17__13__m2s), .qb(),
		.d(n3170), .sdi(n2058), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__13__slave ( .q(_RegFile_17__13), .qb(n2059),
		.d(_RegFile_reg_17__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__14__master ( .q(_RegFile_reg_17__14__m2s), .qb(),
		.d(n3171), .sdi(n2059), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__14__slave ( .q(_RegFile_17__14), .qb(n2060),
		.d(_RegFile_reg_17__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__15__master ( .q(_RegFile_reg_17__15__m2s), .qb(),
		.d(n3172), .sdi(n2060), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__15__slave ( .q(_RegFile_17__15), .qb(n2061),
		.d(_RegFile_reg_17__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__16__master ( .q(_RegFile_reg_17__16__m2s), .qb(),
		.d(n3173), .sdi(n2061), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__16__slave ( .q(_RegFile_17__16), .qb(n2062),
		.d(_RegFile_reg_17__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__17__master ( .q(_RegFile_reg_17__17__m2s), .qb(),
		.d(n3174), .sdi(n2062), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__17__slave ( .q(_RegFile_17__17), .qb(n2063),
		.d(_RegFile_reg_17__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__18__master ( .q(_RegFile_reg_17__18__m2s), .qb(),
		.d(n3175), .sdi(n2063), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__18__slave ( .q(_RegFile_17__18), .qb(n2064),
		.d(_RegFile_reg_17__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__19__master ( .q(_RegFile_reg_17__19__m2s), .qb(),
		.d(n3176), .sdi(n2064), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__19__slave ( .q(_RegFile_17__19), .qb(n2065),
		.d(_RegFile_reg_17__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__1__master ( .q(_RegFile_reg_17__1__m2s), .qb(),
		.d(n3158), .sdi(n4232), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n943),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__1__slave ( .q(_RegFile_17__1), .qb(n4231), .d(_RegFile_reg_17__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n943), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__20__master ( .q(_RegFile_reg_17__20__m2s), .qb(),
		.d(n3177), .sdi(n2065), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__20__slave ( .q(_RegFile_17__20), .qb(n2066),
		.d(_RegFile_reg_17__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__21__master ( .q(_RegFile_reg_17__21__m2s), .qb(),
		.d(n3178), .sdi(n2066), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__21__slave ( .q(_RegFile_17__21), .qb(n2067),
		.d(_RegFile_reg_17__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__22__master ( .q(_RegFile_reg_17__22__m2s), .qb(),
		.d(n3179), .sdi(n2067), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__22__slave ( .q(_RegFile_17__22), .qb(n2068),
		.d(_RegFile_reg_17__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__23__master ( .q(_RegFile_reg_17__23__m2s), .qb(),
		.d(n3180), .sdi(n2068), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__23__slave ( .q(_RegFile_17__23), .qb(n2069),
		.d(_RegFile_reg_17__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__24__master ( .q(_RegFile_reg_17__24__m2s), .qb(),
		.d(n3181), .sdi(n2069), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__24__slave ( .q(_RegFile_17__24), .qb(n2070),
		.d(_RegFile_reg_17__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__25__master ( .q(_RegFile_reg_17__25__m2s), .qb(),
		.d(n3182), .sdi(n2070), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__25__slave ( .q(_RegFile_17__25), .qb(n2071),
		.d(_RegFile_reg_17__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__26__master ( .q(_RegFile_reg_17__26__m2s), .qb(),
		.d(n3183), .sdi(n2071), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__26__slave ( .q(_RegFile_17__26), .qb(n2072),
		.d(_RegFile_reg_17__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__27__master ( .q(_RegFile_reg_17__27__m2s), .qb(),
		.d(n3184), .sdi(n2072), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__27__slave ( .q(_RegFile_17__27), .qb(n2073),
		.d(_RegFile_reg_17__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__28__master ( .q(_RegFile_reg_17__28__m2s), .qb(),
		.d(n3185), .sdi(n2073), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__28__slave ( .q(_RegFile_17__28), .qb(n2074),
		.d(_RegFile_reg_17__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__29__master ( .q(_RegFile_reg_17__29__m2s), .qb(),
		.d(n3186), .sdi(n2074), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__29__slave ( .q(_RegFile_17__29), .qb(n2075),
		.d(_RegFile_reg_17__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__2__master ( .q(_RegFile_reg_17__2__m2s), .qb(),
		.d(n3159), .sdi(n4231), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__2__slave ( .q(_RegFile_17__2), .qb(n4230), .d(_RegFile_reg_17__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__30__master ( .q(_RegFile_reg_17__30__m2s), .qb(),
		.d(n3187), .sdi(n2075), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__30__slave ( .q(_RegFile_17__30), .qb(n2076),
		.d(_RegFile_reg_17__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__31__master ( .q(_RegFile_reg_17__31__m2s), .qb(),
		.d(n3188), .sdi(n2076), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__31__slave ( .q(_RegFile_17__31), .qb(n2077),
		.d(_RegFile_reg_17__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__3__master ( .q(_RegFile_reg_17__3__m2s), .qb(),
		.d(n3160), .sdi(n4230), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__3__slave ( .q(_RegFile_17__3), .qb(n4229), .d(_RegFile_reg_17__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__4__master ( .q(_RegFile_reg_17__4__m2s), .qb(),
		.d(n3161), .sdi(n4229), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__4__slave ( .q(_RegFile_17__4), .qb(n4228), .d(_RegFile_reg_17__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__5__master ( .q(_RegFile_reg_17__5__m2s), .qb(),
		.d(n3162), .sdi(n4228), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__5__slave ( .q(_RegFile_17__5), .qb(n4227), .d(_RegFile_reg_17__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__6__master ( .q(_RegFile_reg_17__6__m2s), .qb(),
		.d(n3163), .sdi(n4227), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__6__slave ( .q(_RegFile_17__6), .qb(n4226), .d(_RegFile_reg_17__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__7__master ( .q(_RegFile_reg_17__7__m2s), .qb(),
		.d(n3164), .sdi(n4226), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__7__slave ( .q(_RegFile_17__7), .qb(n4225), .d(_RegFile_reg_17__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__8__master ( .q(_RegFile_reg_17__8__m2s), .qb(),
		.d(n3165), .sdi(n4225), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__8__slave ( .q(_RegFile_17__8), .qb(n2078), .d(_RegFile_reg_17__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_17__9__master ( .q(_RegFile_reg_17__9__m2s), .qb(),
		.d(n3166), .sdi(n2078), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_17__9__slave ( .q(_RegFile_17__9), .qb(n2079), .d(_RegFile_reg_17__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__0__master ( .q(_RegFile_reg_18__0__m2s), .qb(),
		.d(n3125), .sdi(n2077), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__0__slave ( .q(_RegFile_18__0), .qb(n4224), .d(_RegFile_reg_18__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__10__master ( .q(_RegFile_reg_18__10__m2s), .qb(),
		.d(n3135), .sdi(n2103), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__10__slave ( .q(_RegFile_18__10), .qb(n2080),
		.d(_RegFile_reg_18__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__11__master ( .q(_RegFile_reg_18__11__m2s), .qb(),
		.d(n3136), .sdi(n2080), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__11__slave ( .q(_RegFile_18__11), .qb(n2081),
		.d(_RegFile_reg_18__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__12__master ( .q(_RegFile_reg_18__12__m2s), .qb(),
		.d(n3137), .sdi(n2081), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__12__slave ( .q(_RegFile_18__12), .qb(n2082),
		.d(_RegFile_reg_18__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__13__master ( .q(_RegFile_reg_18__13__m2s), .qb(),
		.d(n3138), .sdi(n2082), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__13__slave ( .q(_RegFile_18__13), .qb(n2083),
		.d(_RegFile_reg_18__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__14__master ( .q(_RegFile_reg_18__14__m2s), .qb(),
		.d(n3139), .sdi(n2083), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__14__slave ( .q(_RegFile_18__14), .qb(n2084),
		.d(_RegFile_reg_18__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__15__master ( .q(_RegFile_reg_18__15__m2s), .qb(),
		.d(n3140), .sdi(n2084), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__15__slave ( .q(_RegFile_18__15), .qb(n2085),
		.d(_RegFile_reg_18__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__16__master ( .q(_RegFile_reg_18__16__m2s), .qb(),
		.d(n3141), .sdi(n2085), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__16__slave ( .q(_RegFile_18__16), .qb(n2086),
		.d(_RegFile_reg_18__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__17__master ( .q(_RegFile_reg_18__17__m2s), .qb(),
		.d(n3142), .sdi(n2086), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__17__slave ( .q(_RegFile_18__17), .qb(n2087),
		.d(_RegFile_reg_18__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__18__master ( .q(_RegFile_reg_18__18__m2s), .qb(),
		.d(n3143), .sdi(n2087), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__18__slave ( .q(_RegFile_18__18), .qb(n2088),
		.d(_RegFile_reg_18__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__19__master ( .q(_RegFile_reg_18__19__m2s), .qb(),
		.d(n3144), .sdi(n2088), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__19__slave ( .q(_RegFile_18__19), .qb(n2089),
		.d(_RegFile_reg_18__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__1__master ( .q(_RegFile_reg_18__1__m2s), .qb(),
		.d(n3126), .sdi(n4224), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n942),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__1__slave ( .q(_RegFile_18__1), .qb(n4223), .d(_RegFile_reg_18__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n942), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__20__master ( .q(_RegFile_reg_18__20__m2s), .qb(),
		.d(n3145), .sdi(n2089), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__20__slave ( .q(_RegFile_18__20), .qb(n2090),
		.d(_RegFile_reg_18__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__21__master ( .q(_RegFile_reg_18__21__m2s), .qb(),
		.d(n3146), .sdi(n2090), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__21__slave ( .q(_RegFile_18__21), .qb(n2091),
		.d(_RegFile_reg_18__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__22__master ( .q(_RegFile_reg_18__22__m2s), .qb(),
		.d(n3147), .sdi(n2091), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__22__slave ( .q(_RegFile_18__22), .qb(n2092),
		.d(_RegFile_reg_18__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__23__master ( .q(_RegFile_reg_18__23__m2s), .qb(),
		.d(n3148), .sdi(n2092), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__23__slave ( .q(_RegFile_18__23), .qb(n2093),
		.d(_RegFile_reg_18__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__24__master ( .q(_RegFile_reg_18__24__m2s), .qb(),
		.d(n3149), .sdi(n2093), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__24__slave ( .q(_RegFile_18__24), .qb(n2094),
		.d(_RegFile_reg_18__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__25__master ( .q(_RegFile_reg_18__25__m2s), .qb(),
		.d(n3150), .sdi(n2094), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__25__slave ( .q(_RegFile_18__25), .qb(n2095),
		.d(_RegFile_reg_18__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__26__master ( .q(_RegFile_reg_18__26__m2s), .qb(),
		.d(n3151), .sdi(n2095), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__26__slave ( .q(_RegFile_18__26), .qb(n2096),
		.d(_RegFile_reg_18__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__27__master ( .q(_RegFile_reg_18__27__m2s), .qb(),
		.d(n3152), .sdi(n2096), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__27__slave ( .q(_RegFile_18__27), .qb(n2097),
		.d(_RegFile_reg_18__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__28__master ( .q(_RegFile_reg_18__28__m2s), .qb(),
		.d(n3153), .sdi(n2097), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__28__slave ( .q(_RegFile_18__28), .qb(n2098),
		.d(_RegFile_reg_18__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__29__master ( .q(_RegFile_reg_18__29__m2s), .qb(),
		.d(n3154), .sdi(n2098), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__29__slave ( .q(_RegFile_18__29), .qb(n2099),
		.d(_RegFile_reg_18__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__2__master ( .q(_RegFile_reg_18__2__m2s), .qb(),
		.d(n3127), .sdi(n4223), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n961),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__2__slave ( .q(_RegFile_18__2), .qb(n4222), .d(_RegFile_reg_18__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n961), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__30__master ( .q(_RegFile_reg_18__30__m2s), .qb(),
		.d(n3155), .sdi(n2099), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__30__slave ( .q(_RegFile_18__30), .qb(n2100),
		.d(_RegFile_reg_18__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__31__master ( .q(_RegFile_reg_18__31__m2s), .qb(),
		.d(n3156), .sdi(n2100), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__31__slave ( .q(_RegFile_18__31), .qb(n2101),
		.d(_RegFile_reg_18__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__3__master ( .q(_RegFile_reg_18__3__m2s), .qb(),
		.d(n3128), .sdi(n4222), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__3__slave ( .q(_RegFile_18__3), .qb(n4221), .d(_RegFile_reg_18__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__4__master ( .q(_RegFile_reg_18__4__m2s), .qb(),
		.d(n3129), .sdi(n4221), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__4__slave ( .q(_RegFile_18__4), .qb(n4220), .d(_RegFile_reg_18__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__5__master ( .q(_RegFile_reg_18__5__m2s), .qb(),
		.d(n3130), .sdi(n4220), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__5__slave ( .q(_RegFile_18__5), .qb(n4219), .d(_RegFile_reg_18__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__6__master ( .q(_RegFile_reg_18__6__m2s), .qb(),
		.d(n3131), .sdi(n4219), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__6__slave ( .q(_RegFile_18__6), .qb(n4218), .d(_RegFile_reg_18__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__7__master ( .q(_RegFile_reg_18__7__m2s), .qb(),
		.d(n3132), .sdi(n4218), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__7__slave ( .q(_RegFile_18__7), .qb(n4217), .d(_RegFile_reg_18__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__8__master ( .q(_RegFile_reg_18__8__m2s), .qb(),
		.d(n3133), .sdi(n4217), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__8__slave ( .q(_RegFile_18__8), .qb(n2102), .d(_RegFile_reg_18__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_18__9__master ( .q(_RegFile_reg_18__9__m2s), .qb(),
		.d(n3134), .sdi(n2102), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_18__9__slave ( .q(_RegFile_18__9), .qb(n2103), .d(_RegFile_reg_18__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__0__master ( .q(_RegFile_reg_19__0__m2s), .qb(),
		.d(n3093), .sdi(n2101), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__0__slave ( .q(_RegFile_19__0), .qb(n4216), .d(_RegFile_reg_19__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__10__master ( .q(_RegFile_reg_19__10__m2s), .qb(),
		.d(n3103), .sdi(n2127), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__10__slave ( .q(_RegFile_19__10), .qb(n2104),
		.d(_RegFile_reg_19__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__11__master ( .q(_RegFile_reg_19__11__m2s), .qb(),
		.d(n3104), .sdi(n2104), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__11__slave ( .q(_RegFile_19__11), .qb(n2105),
		.d(_RegFile_reg_19__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__12__master ( .q(_RegFile_reg_19__12__m2s), .qb(),
		.d(n3105), .sdi(n2105), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__12__slave ( .q(_RegFile_19__12), .qb(n2106),
		.d(_RegFile_reg_19__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__13__master ( .q(_RegFile_reg_19__13__m2s), .qb(),
		.d(n3106), .sdi(n2106), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__13__slave ( .q(_RegFile_19__13), .qb(n2107),
		.d(_RegFile_reg_19__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__14__master ( .q(_RegFile_reg_19__14__m2s), .qb(),
		.d(n3107), .sdi(n2107), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__14__slave ( .q(_RegFile_19__14), .qb(n2108),
		.d(_RegFile_reg_19__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__15__master ( .q(_RegFile_reg_19__15__m2s), .qb(),
		.d(n3108), .sdi(n2108), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__15__slave ( .q(_RegFile_19__15), .qb(n2109),
		.d(_RegFile_reg_19__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__16__master ( .q(_RegFile_reg_19__16__m2s), .qb(),
		.d(n3109), .sdi(n2109), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__16__slave ( .q(_RegFile_19__16), .qb(n2110),
		.d(_RegFile_reg_19__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__17__master ( .q(_RegFile_reg_19__17__m2s), .qb(),
		.d(n3110), .sdi(n2110), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__17__slave ( .q(_RegFile_19__17), .qb(n2111),
		.d(_RegFile_reg_19__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__18__master ( .q(_RegFile_reg_19__18__m2s), .qb(),
		.d(n3111), .sdi(n2111), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__18__slave ( .q(_RegFile_19__18), .qb(n2112),
		.d(_RegFile_reg_19__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__19__master ( .q(_RegFile_reg_19__19__m2s), .qb(),
		.d(n3112), .sdi(n2112), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__19__slave ( .q(_RegFile_19__19), .qb(n2113),
		.d(_RegFile_reg_19__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__1__master ( .q(_RegFile_reg_19__1__m2s), .qb(),
		.d(n3094), .sdi(n4216), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n941),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__1__slave ( .q(_RegFile_19__1), .qb(n4215), .d(_RegFile_reg_19__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n941), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__20__master ( .q(_RegFile_reg_19__20__m2s), .qb(),
		.d(n3113), .sdi(n2113), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__20__slave ( .q(_RegFile_19__20), .qb(n2114),
		.d(_RegFile_reg_19__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__21__master ( .q(_RegFile_reg_19__21__m2s), .qb(),
		.d(n3114), .sdi(n2114), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__21__slave ( .q(_RegFile_19__21), .qb(n2115),
		.d(_RegFile_reg_19__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__22__master ( .q(_RegFile_reg_19__22__m2s), .qb(),
		.d(n3115), .sdi(n2115), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__22__slave ( .q(_RegFile_19__22), .qb(n2116),
		.d(_RegFile_reg_19__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__23__master ( .q(_RegFile_reg_19__23__m2s), .qb(),
		.d(n3116), .sdi(n2116), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__23__slave ( .q(_RegFile_19__23), .qb(n2117),
		.d(_RegFile_reg_19__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__24__master ( .q(_RegFile_reg_19__24__m2s), .qb(),
		.d(n3117), .sdi(n2117), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__24__slave ( .q(_RegFile_19__24), .qb(n2118),
		.d(_RegFile_reg_19__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__25__master ( .q(_RegFile_reg_19__25__m2s), .qb(),
		.d(n3118), .sdi(n2118), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__25__slave ( .q(_RegFile_19__25), .qb(n2119),
		.d(_RegFile_reg_19__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__26__master ( .q(_RegFile_reg_19__26__m2s), .qb(),
		.d(n3119), .sdi(n2119), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__26__slave ( .q(_RegFile_19__26), .qb(n2120),
		.d(_RegFile_reg_19__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__27__master ( .q(_RegFile_reg_19__27__m2s), .qb(),
		.d(n3120), .sdi(n2120), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__27__slave ( .q(_RegFile_19__27), .qb(n2121),
		.d(_RegFile_reg_19__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__28__master ( .q(_RegFile_reg_19__28__m2s), .qb(),
		.d(n3121), .sdi(n2121), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__28__slave ( .q(_RegFile_19__28), .qb(n2122),
		.d(_RegFile_reg_19__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__29__master ( .q(_RegFile_reg_19__29__m2s), .qb(),
		.d(n3122), .sdi(n2122), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__29__slave ( .q(_RegFile_19__29), .qb(n2123),
		.d(_RegFile_reg_19__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__2__master ( .q(_RegFile_reg_19__2__m2s), .qb(),
		.d(n3095), .sdi(n4215), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__2__slave ( .q(_RegFile_19__2), .qb(n4214), .d(_RegFile_reg_19__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__30__master ( .q(_RegFile_reg_19__30__m2s), .qb(),
		.d(n3123), .sdi(n2123), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__30__slave ( .q(_RegFile_19__30), .qb(n2124),
		.d(_RegFile_reg_19__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__31__master ( .q(_RegFile_reg_19__31__m2s), .qb(),
		.d(n3124), .sdi(n2124), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__31__slave ( .q(_RegFile_19__31), .qb(n2125),
		.d(_RegFile_reg_19__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__3__master ( .q(_RegFile_reg_19__3__m2s), .qb(),
		.d(n3096), .sdi(n4214), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__3__slave ( .q(_RegFile_19__3), .qb(n4213), .d(_RegFile_reg_19__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__4__master ( .q(_RegFile_reg_19__4__m2s), .qb(),
		.d(n3097), .sdi(n4213), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__4__slave ( .q(_RegFile_19__4), .qb(n4212), .d(_RegFile_reg_19__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__5__master ( .q(_RegFile_reg_19__5__m2s), .qb(),
		.d(n3098), .sdi(n4212), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__5__slave ( .q(_RegFile_19__5), .qb(n4211), .d(_RegFile_reg_19__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__6__master ( .q(_RegFile_reg_19__6__m2s), .qb(),
		.d(n3099), .sdi(n4211), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__6__slave ( .q(_RegFile_19__6), .qb(n4210), .d(_RegFile_reg_19__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__7__master ( .q(_RegFile_reg_19__7__m2s), .qb(),
		.d(n3100), .sdi(n4210), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__7__slave ( .q(_RegFile_19__7), .qb(n4209), .d(_RegFile_reg_19__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__8__master ( .q(_RegFile_reg_19__8__m2s), .qb(),
		.d(n3101), .sdi(n4209), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__8__slave ( .q(_RegFile_19__8), .qb(n2126), .d(_RegFile_reg_19__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_19__9__master ( .q(_RegFile_reg_19__9__m2s), .qb(),
		.d(n3102), .sdi(n2126), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n940),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_19__9__slave ( .q(_RegFile_19__9), .qb(n2127), .d(_RegFile_reg_19__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n940), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__0__master ( .q(_RegFile_reg_1__0__m2s), .qb(),
		.d(n3669), .sdi(n1885), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__0__slave ( .q(_RegFile_1__0), .qb(n4360), .d(_RegFile_reg_1__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__10__master ( .q(_RegFile_reg_1__10__m2s), .qb(),
		.d(n3679), .sdi(n2151), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__10__slave ( .q(_RegFile_1__10), .qb(n2128), .d(_RegFile_reg_1__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__11__master ( .q(_RegFile_reg_1__11__m2s), .qb(),
		.d(n3680), .sdi(n2128), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__11__slave ( .q(_RegFile_1__11), .qb(n2129), .d(_RegFile_reg_1__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__12__master ( .q(_RegFile_reg_1__12__m2s), .qb(),
		.d(n3681), .sdi(n2129), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__12__slave ( .q(_RegFile_1__12), .qb(n2130), .d(_RegFile_reg_1__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__13__master ( .q(_RegFile_reg_1__13__m2s), .qb(),
		.d(n3682), .sdi(n2130), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__13__slave ( .q(_RegFile_1__13), .qb(n2131), .d(_RegFile_reg_1__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__14__master ( .q(_RegFile_reg_1__14__m2s), .qb(),
		.d(n3683), .sdi(n2131), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__14__slave ( .q(_RegFile_1__14), .qb(n2132), .d(_RegFile_reg_1__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__15__master ( .q(_RegFile_reg_1__15__m2s), .qb(),
		.d(n3684), .sdi(n2132), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__15__slave ( .q(_RegFile_1__15), .qb(n2133), .d(_RegFile_reg_1__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__16__master ( .q(_RegFile_reg_1__16__m2s), .qb(),
		.d(n3685), .sdi(n2133), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__16__slave ( .q(_RegFile_1__16), .qb(n2134), .d(_RegFile_reg_1__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__17__master ( .q(_RegFile_reg_1__17__m2s), .qb(),
		.d(n3686), .sdi(n2134), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__17__slave ( .q(_RegFile_1__17), .qb(n2135), .d(_RegFile_reg_1__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__18__master ( .q(_RegFile_reg_1__18__m2s), .qb(),
		.d(n3687), .sdi(n2135), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__18__slave ( .q(_RegFile_1__18), .qb(n2136), .d(_RegFile_reg_1__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__19__master ( .q(_RegFile_reg_1__19__m2s), .qb(),
		.d(n3688), .sdi(n2136), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__19__slave ( .q(_RegFile_1__19), .qb(n2137), .d(_RegFile_reg_1__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__1__master ( .q(_RegFile_reg_1__1__m2s), .qb(),
		.d(n3670), .sdi(n4360), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__1__slave ( .q(_RegFile_1__1), .qb(n4359), .d(_RegFile_reg_1__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__20__master ( .q(_RegFile_reg_1__20__m2s), .qb(),
		.d(n3689), .sdi(n2137), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__20__slave ( .q(_RegFile_1__20), .qb(n2138), .d(_RegFile_reg_1__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__21__master ( .q(_RegFile_reg_1__21__m2s), .qb(),
		.d(n3690), .sdi(n2138), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__21__slave ( .q(_RegFile_1__21), .qb(n2139), .d(_RegFile_reg_1__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__22__master ( .q(_RegFile_reg_1__22__m2s), .qb(),
		.d(n3691), .sdi(n2139), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__22__slave ( .q(_RegFile_1__22), .qb(n2140), .d(_RegFile_reg_1__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__23__master ( .q(_RegFile_reg_1__23__m2s), .qb(),
		.d(n3692), .sdi(n2140), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__23__slave ( .q(_RegFile_1__23), .qb(n2141), .d(_RegFile_reg_1__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__24__master ( .q(_RegFile_reg_1__24__m2s), .qb(),
		.d(n3693), .sdi(n2141), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__24__slave ( .q(_RegFile_1__24), .qb(n2142), .d(_RegFile_reg_1__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__25__master ( .q(_RegFile_reg_1__25__m2s), .qb(),
		.d(n3694), .sdi(n2142), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__25__slave ( .q(_RegFile_1__25), .qb(n2143), .d(_RegFile_reg_1__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__26__master ( .q(_RegFile_reg_1__26__m2s), .qb(),
		.d(n3695), .sdi(n2143), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__26__slave ( .q(_RegFile_1__26), .qb(n2144), .d(_RegFile_reg_1__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__27__master ( .q(_RegFile_reg_1__27__m2s), .qb(),
		.d(n3696), .sdi(n2144), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__27__slave ( .q(_RegFile_1__27), .qb(n2145), .d(_RegFile_reg_1__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__28__master ( .q(_RegFile_reg_1__28__m2s), .qb(),
		.d(n3697), .sdi(n2145), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__28__slave ( .q(_RegFile_1__28), .qb(n2146), .d(_RegFile_reg_1__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__29__master ( .q(_RegFile_reg_1__29__m2s), .qb(),
		.d(n3698), .sdi(n2146), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__29__slave ( .q(_RegFile_1__29), .qb(n2147), .d(_RegFile_reg_1__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__2__master ( .q(_RegFile_reg_1__2__m2s), .qb(),
		.d(n3671), .sdi(n4359), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n962),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__2__slave ( .q(_RegFile_1__2), .qb(n4358), .d(_RegFile_reg_1__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n962), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__30__master ( .q(_RegFile_reg_1__30__m2s), .qb(),
		.d(n3699), .sdi(n2147), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__30__slave ( .q(_RegFile_1__30), .qb(n2148), .d(_RegFile_reg_1__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__31__master ( .q(_RegFile_reg_1__31__m2s), .qb(),
		.d(n3700), .sdi(n2148), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__31__slave ( .q(_RegFile_1__31), .qb(n2149), .d(_RegFile_reg_1__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__3__master ( .q(_RegFile_reg_1__3__m2s), .qb(),
		.d(n3672), .sdi(n4358), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__3__slave ( .q(_RegFile_1__3), .qb(n4357), .d(_RegFile_reg_1__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__4__master ( .q(_RegFile_reg_1__4__m2s), .qb(),
		.d(n3673), .sdi(n4357), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__4__slave ( .q(_RegFile_1__4), .qb(n4356), .d(_RegFile_reg_1__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__5__master ( .q(_RegFile_reg_1__5__m2s), .qb(),
		.d(n3674), .sdi(n4356), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__5__slave ( .q(_RegFile_1__5), .qb(n4355), .d(_RegFile_reg_1__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__6__master ( .q(_RegFile_reg_1__6__m2s), .qb(),
		.d(n3675), .sdi(n4355), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__6__slave ( .q(_RegFile_1__6), .qb(n4354), .d(_RegFile_reg_1__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__7__master ( .q(_RegFile_reg_1__7__m2s), .qb(),
		.d(n3676), .sdi(n4354), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n939),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__7__slave ( .q(_RegFile_1__7), .qb(n4353), .d(_RegFile_reg_1__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n939), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__8__master ( .q(_RegFile_reg_1__8__m2s), .qb(),
		.d(n3677), .sdi(n4353), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__8__slave ( .q(_RegFile_1__8), .qb(n2150), .d(_RegFile_reg_1__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_1__9__master ( .q(_RegFile_reg_1__9__m2s), .qb(),
		.d(n3678), .sdi(n2150), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_1__9__slave ( .q(_RegFile_1__9), .qb(n2151), .d(_RegFile_reg_1__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__0__master ( .q(_RegFile_reg_20__0__m2s), .qb(),
		.d(n3061), .sdi(n2125), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__0__slave ( .q(_RegFile_20__0), .qb(n4208), .d(_RegFile_reg_20__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__10__master ( .q(_RegFile_reg_20__10__m2s), .qb(),
		.d(n3071), .sdi(n2175), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__10__slave ( .q(_RegFile_20__10), .qb(n2152),
		.d(_RegFile_reg_20__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__11__master ( .q(_RegFile_reg_20__11__m2s), .qb(),
		.d(n3072), .sdi(n2152), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__11__slave ( .q(_RegFile_20__11), .qb(n2153),
		.d(_RegFile_reg_20__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__12__master ( .q(_RegFile_reg_20__12__m2s), .qb(),
		.d(n3073), .sdi(n2153), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__12__slave ( .q(_RegFile_20__12), .qb(n2154),
		.d(_RegFile_reg_20__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__13__master ( .q(_RegFile_reg_20__13__m2s), .qb(),
		.d(n3074), .sdi(n2154), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__13__slave ( .q(_RegFile_20__13), .qb(n2155),
		.d(_RegFile_reg_20__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__14__master ( .q(_RegFile_reg_20__14__m2s), .qb(),
		.d(n3075), .sdi(n2155), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__14__slave ( .q(_RegFile_20__14), .qb(n2156),
		.d(_RegFile_reg_20__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__15__master ( .q(_RegFile_reg_20__15__m2s), .qb(),
		.d(n3076), .sdi(n2156), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__15__slave ( .q(_RegFile_20__15), .qb(n2157),
		.d(_RegFile_reg_20__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__16__master ( .q(_RegFile_reg_20__16__m2s), .qb(),
		.d(n3077), .sdi(n2157), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__16__slave ( .q(_RegFile_20__16), .qb(n2158),
		.d(_RegFile_reg_20__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__17__master ( .q(_RegFile_reg_20__17__m2s), .qb(),
		.d(n3078), .sdi(n2158), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__17__slave ( .q(_RegFile_20__17), .qb(n2159),
		.d(_RegFile_reg_20__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__18__master ( .q(_RegFile_reg_20__18__m2s), .qb(),
		.d(n3079), .sdi(n2159), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__18__slave ( .q(_RegFile_20__18), .qb(n2160),
		.d(_RegFile_reg_20__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__19__master ( .q(_RegFile_reg_20__19__m2s), .qb(),
		.d(n3080), .sdi(n2160), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__19__slave ( .q(_RegFile_20__19), .qb(n2161),
		.d(_RegFile_reg_20__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__1__master ( .q(_RegFile_reg_20__1__m2s), .qb(),
		.d(n3062), .sdi(n4208), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__1__slave ( .q(_RegFile_20__1), .qb(n4207), .d(_RegFile_reg_20__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__20__master ( .q(_RegFile_reg_20__20__m2s), .qb(),
		.d(n3081), .sdi(n2161), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__20__slave ( .q(_RegFile_20__20), .qb(n2162),
		.d(_RegFile_reg_20__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__21__master ( .q(_RegFile_reg_20__21__m2s), .qb(),
		.d(n3082), .sdi(n2162), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__21__slave ( .q(_RegFile_20__21), .qb(n2163),
		.d(_RegFile_reg_20__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__22__master ( .q(_RegFile_reg_20__22__m2s), .qb(),
		.d(n3083), .sdi(n2163), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__22__slave ( .q(_RegFile_20__22), .qb(n2164),
		.d(_RegFile_reg_20__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__23__master ( .q(_RegFile_reg_20__23__m2s), .qb(),
		.d(n3084), .sdi(n2164), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__23__slave ( .q(_RegFile_20__23), .qb(n2165),
		.d(_RegFile_reg_20__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__24__master ( .q(_RegFile_reg_20__24__m2s), .qb(),
		.d(n3085), .sdi(n2165), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__24__slave ( .q(_RegFile_20__24), .qb(n2166),
		.d(_RegFile_reg_20__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__25__master ( .q(_RegFile_reg_20__25__m2s), .qb(),
		.d(n3086), .sdi(n2166), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__25__slave ( .q(_RegFile_20__25), .qb(n2167),
		.d(_RegFile_reg_20__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__26__master ( .q(_RegFile_reg_20__26__m2s), .qb(),
		.d(n3087), .sdi(n2167), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__26__slave ( .q(_RegFile_20__26), .qb(n2168),
		.d(_RegFile_reg_20__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__27__master ( .q(_RegFile_reg_20__27__m2s), .qb(),
		.d(n3088), .sdi(n2168), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__27__slave ( .q(_RegFile_20__27), .qb(n2169),
		.d(_RegFile_reg_20__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__28__master ( .q(_RegFile_reg_20__28__m2s), .qb(),
		.d(n3089), .sdi(n2169), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__28__slave ( .q(_RegFile_20__28), .qb(n2170),
		.d(_RegFile_reg_20__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__29__master ( .q(_RegFile_reg_20__29__m2s), .qb(),
		.d(n3090), .sdi(n2170), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__29__slave ( .q(_RegFile_20__29), .qb(n2171),
		.d(_RegFile_reg_20__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__2__master ( .q(_RegFile_reg_20__2__m2s), .qb(),
		.d(n3063), .sdi(n4207), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n963),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__2__slave ( .q(_RegFile_20__2), .qb(n4206), .d(_RegFile_reg_20__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n963), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__30__master ( .q(_RegFile_reg_20__30__m2s), .qb(),
		.d(n3091), .sdi(n2171), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__30__slave ( .q(_RegFile_20__30), .qb(n2172),
		.d(_RegFile_reg_20__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__31__master ( .q(_RegFile_reg_20__31__m2s), .qb(),
		.d(n3092), .sdi(n2172), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__31__slave ( .q(_RegFile_20__31), .qb(n2173),
		.d(_RegFile_reg_20__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__3__master ( .q(_RegFile_reg_20__3__m2s), .qb(),
		.d(n3064), .sdi(n4206), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__3__slave ( .q(_RegFile_20__3), .qb(n4205), .d(_RegFile_reg_20__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__4__master ( .q(_RegFile_reg_20__4__m2s), .qb(),
		.d(n3065), .sdi(n4205), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__4__slave ( .q(_RegFile_20__4), .qb(n4204), .d(_RegFile_reg_20__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__5__master ( .q(_RegFile_reg_20__5__m2s), .qb(),
		.d(n3066), .sdi(n4204), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__5__slave ( .q(_RegFile_20__5), .qb(n4203), .d(_RegFile_reg_20__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__6__master ( .q(_RegFile_reg_20__6__m2s), .qb(),
		.d(n3067), .sdi(n4203), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__6__slave ( .q(_RegFile_20__6), .qb(n4202), .d(_RegFile_reg_20__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__7__master ( .q(_RegFile_reg_20__7__m2s), .qb(),
		.d(n3068), .sdi(n4202), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__7__slave ( .q(_RegFile_20__7), .qb(n4201), .d(_RegFile_reg_20__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__8__master ( .q(_RegFile_reg_20__8__m2s), .qb(),
		.d(n3069), .sdi(n4201), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__8__slave ( .q(_RegFile_20__8), .qb(n2174), .d(_RegFile_reg_20__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_20__9__master ( .q(_RegFile_reg_20__9__m2s), .qb(),
		.d(n3070), .sdi(n2174), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_20__9__slave ( .q(_RegFile_20__9), .qb(n2175), .d(_RegFile_reg_20__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__0__master ( .q(_RegFile_reg_21__0__m2s), .qb(),
		.d(n3029), .sdi(n2173), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__0__slave ( .q(_RegFile_21__0), .qb(n4200), .d(_RegFile_reg_21__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__10__master ( .q(_RegFile_reg_21__10__m2s), .qb(),
		.d(n3039), .sdi(n2199), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__10__slave ( .q(_RegFile_21__10), .qb(n2176),
		.d(_RegFile_reg_21__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__11__master ( .q(_RegFile_reg_21__11__m2s), .qb(),
		.d(n3040), .sdi(n2176), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__11__slave ( .q(_RegFile_21__11), .qb(n2177),
		.d(_RegFile_reg_21__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__12__master ( .q(_RegFile_reg_21__12__m2s), .qb(),
		.d(n3041), .sdi(n2177), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__12__slave ( .q(_RegFile_21__12), .qb(n2178),
		.d(_RegFile_reg_21__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__13__master ( .q(_RegFile_reg_21__13__m2s), .qb(),
		.d(n3042), .sdi(n2178), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__13__slave ( .q(_RegFile_21__13), .qb(n2179),
		.d(_RegFile_reg_21__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__14__master ( .q(_RegFile_reg_21__14__m2s), .qb(),
		.d(n3043), .sdi(n2179), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__14__slave ( .q(_RegFile_21__14), .qb(n2180),
		.d(_RegFile_reg_21__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__15__master ( .q(_RegFile_reg_21__15__m2s), .qb(),
		.d(n3044), .sdi(n2180), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__15__slave ( .q(_RegFile_21__15), .qb(n2181),
		.d(_RegFile_reg_21__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__16__master ( .q(_RegFile_reg_21__16__m2s), .qb(),
		.d(n3045), .sdi(n2181), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__16__slave ( .q(_RegFile_21__16), .qb(n2182),
		.d(_RegFile_reg_21__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__17__master ( .q(_RegFile_reg_21__17__m2s), .qb(),
		.d(n3046), .sdi(n2182), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__17__slave ( .q(_RegFile_21__17), .qb(n2183),
		.d(_RegFile_reg_21__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__18__master ( .q(_RegFile_reg_21__18__m2s), .qb(),
		.d(n3047), .sdi(n2183), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n964),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__18__slave ( .q(_RegFile_21__18), .qb(n2184),
		.d(_RegFile_reg_21__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n964), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__19__master ( .q(_RegFile_reg_21__19__m2s), .qb(),
		.d(n3048), .sdi(n2184), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__19__slave ( .q(_RegFile_21__19), .qb(n2185),
		.d(_RegFile_reg_21__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__1__master ( .q(_RegFile_reg_21__1__m2s), .qb(),
		.d(n3030), .sdi(n4200), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__1__slave ( .q(_RegFile_21__1), .qb(n4199), .d(_RegFile_reg_21__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__20__master ( .q(_RegFile_reg_21__20__m2s), .qb(),
		.d(n3049), .sdi(n2185), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__20__slave ( .q(_RegFile_21__20), .qb(n2186),
		.d(_RegFile_reg_21__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__21__master ( .q(_RegFile_reg_21__21__m2s), .qb(),
		.d(n3050), .sdi(n2186), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__21__slave ( .q(_RegFile_21__21), .qb(n2187),
		.d(_RegFile_reg_21__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__22__master ( .q(_RegFile_reg_21__22__m2s), .qb(),
		.d(n3051), .sdi(n2187), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__22__slave ( .q(_RegFile_21__22), .qb(n2188),
		.d(_RegFile_reg_21__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__23__master ( .q(_RegFile_reg_21__23__m2s), .qb(),
		.d(n3052), .sdi(n2188), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__23__slave ( .q(_RegFile_21__23), .qb(n2189),
		.d(_RegFile_reg_21__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__24__master ( .q(_RegFile_reg_21__24__m2s), .qb(),
		.d(n3053), .sdi(n2189), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__24__slave ( .q(_RegFile_21__24), .qb(n2190),
		.d(_RegFile_reg_21__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__25__master ( .q(_RegFile_reg_21__25__m2s), .qb(),
		.d(n3054), .sdi(n2190), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__25__slave ( .q(_RegFile_21__25), .qb(n2191),
		.d(_RegFile_reg_21__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__26__master ( .q(_RegFile_reg_21__26__m2s), .qb(),
		.d(n3055), .sdi(n2191), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__26__slave ( .q(_RegFile_21__26), .qb(n2192),
		.d(_RegFile_reg_21__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__27__master ( .q(_RegFile_reg_21__27__m2s), .qb(),
		.d(n3056), .sdi(n2192), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__27__slave ( .q(_RegFile_21__27), .qb(n2193),
		.d(_RegFile_reg_21__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__28__master ( .q(_RegFile_reg_21__28__m2s), .qb(),
		.d(n3057), .sdi(n2193), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__28__slave ( .q(_RegFile_21__28), .qb(n2194),
		.d(_RegFile_reg_21__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__29__master ( .q(_RegFile_reg_21__29__m2s), .qb(),
		.d(n3058), .sdi(n2194), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__29__slave ( .q(_RegFile_21__29), .qb(n2195),
		.d(_RegFile_reg_21__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__2__master ( .q(_RegFile_reg_21__2__m2s), .qb(),
		.d(n3031), .sdi(n4199), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__2__slave ( .q(_RegFile_21__2), .qb(n4198), .d(_RegFile_reg_21__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__30__master ( .q(_RegFile_reg_21__30__m2s), .qb(),
		.d(n3059), .sdi(n2195), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__30__slave ( .q(_RegFile_21__30), .qb(n2196),
		.d(_RegFile_reg_21__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__31__master ( .q(_RegFile_reg_21__31__m2s), .qb(),
		.d(n3060), .sdi(n2196), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__31__slave ( .q(_RegFile_21__31), .qb(n2197),
		.d(_RegFile_reg_21__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__3__master ( .q(_RegFile_reg_21__3__m2s), .qb(),
		.d(n3032), .sdi(n4198), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n937),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__3__slave ( .q(_RegFile_21__3), .qb(n4197), .d(_RegFile_reg_21__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n937), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__4__master ( .q(_RegFile_reg_21__4__m2s), .qb(),
		.d(n3033), .sdi(n4197), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__4__slave ( .q(_RegFile_21__4), .qb(n4196), .d(_RegFile_reg_21__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__5__master ( .q(_RegFile_reg_21__5__m2s), .qb(),
		.d(n3034), .sdi(n4196), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__5__slave ( .q(_RegFile_21__5), .qb(n4195), .d(_RegFile_reg_21__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__6__master ( .q(_RegFile_reg_21__6__m2s), .qb(),
		.d(n3035), .sdi(n4195), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__6__slave ( .q(_RegFile_21__6), .qb(n4194), .d(_RegFile_reg_21__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__7__master ( .q(_RegFile_reg_21__7__m2s), .qb(),
		.d(n3036), .sdi(n4194), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__7__slave ( .q(_RegFile_21__7), .qb(n4193), .d(_RegFile_reg_21__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__8__master ( .q(_RegFile_reg_21__8__m2s), .qb(),
		.d(n3037), .sdi(n4193), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__8__slave ( .q(_RegFile_21__8), .qb(n2198), .d(_RegFile_reg_21__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_21__9__master ( .q(_RegFile_reg_21__9__m2s), .qb(),
		.d(n3038), .sdi(n2198), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_21__9__slave ( .q(_RegFile_21__9), .qb(n2199), .d(_RegFile_reg_21__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__0__master ( .q(_RegFile_reg_22__0__m2s), .qb(),
		.d(n2997), .sdi(n2197), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__0__slave ( .q(_RegFile_22__0), .qb(n4192), .d(_RegFile_reg_22__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__10__master ( .q(_RegFile_reg_22__10__m2s), .qb(),
		.d(n3007), .sdi(n2223), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__10__slave ( .q(_RegFile_22__10), .qb(n2200),
		.d(_RegFile_reg_22__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__11__master ( .q(_RegFile_reg_22__11__m2s), .qb(),
		.d(n3008), .sdi(n2200), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__11__slave ( .q(_RegFile_22__11), .qb(n2201),
		.d(_RegFile_reg_22__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__12__master ( .q(_RegFile_reg_22__12__m2s), .qb(),
		.d(n3009), .sdi(n2201), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__12__slave ( .q(_RegFile_22__12), .qb(n2202),
		.d(_RegFile_reg_22__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__13__master ( .q(_RegFile_reg_22__13__m2s), .qb(),
		.d(n3010), .sdi(n2202), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__13__slave ( .q(_RegFile_22__13), .qb(n2203),
		.d(_RegFile_reg_22__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__14__master ( .q(_RegFile_reg_22__14__m2s), .qb(),
		.d(n3011), .sdi(n2203), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__14__slave ( .q(_RegFile_22__14), .qb(n2204),
		.d(_RegFile_reg_22__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__15__master ( .q(_RegFile_reg_22__15__m2s), .qb(),
		.d(n3012), .sdi(n2204), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__15__slave ( .q(_RegFile_22__15), .qb(n2205),
		.d(_RegFile_reg_22__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__16__master ( .q(_RegFile_reg_22__16__m2s), .qb(),
		.d(n3013), .sdi(n2205), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n965),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__16__slave ( .q(_RegFile_22__16), .qb(n2206),
		.d(_RegFile_reg_22__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n965), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__17__master ( .q(_RegFile_reg_22__17__m2s), .qb(),
		.d(n3014), .sdi(n2206), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__17__slave ( .q(_RegFile_22__17), .qb(n2207),
		.d(_RegFile_reg_22__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__18__master ( .q(_RegFile_reg_22__18__m2s), .qb(),
		.d(n3015), .sdi(n2207), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__18__slave ( .q(_RegFile_22__18), .qb(n2208),
		.d(_RegFile_reg_22__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__19__master ( .q(_RegFile_reg_22__19__m2s), .qb(),
		.d(n3016), .sdi(n2208), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__19__slave ( .q(_RegFile_22__19), .qb(n2209),
		.d(_RegFile_reg_22__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__1__master ( .q(_RegFile_reg_22__1__m2s), .qb(),
		.d(n2998), .sdi(n4192), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__1__slave ( .q(_RegFile_22__1), .qb(n4191), .d(_RegFile_reg_22__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__20__master ( .q(_RegFile_reg_22__20__m2s), .qb(),
		.d(n3017), .sdi(n2209), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__20__slave ( .q(_RegFile_22__20), .qb(n2210),
		.d(_RegFile_reg_22__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__21__master ( .q(_RegFile_reg_22__21__m2s), .qb(),
		.d(n3018), .sdi(n2210), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__21__slave ( .q(_RegFile_22__21), .qb(n2211),
		.d(_RegFile_reg_22__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__22__master ( .q(_RegFile_reg_22__22__m2s), .qb(),
		.d(n3019), .sdi(n2211), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__22__slave ( .q(_RegFile_22__22), .qb(n2212),
		.d(_RegFile_reg_22__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__23__master ( .q(_RegFile_reg_22__23__m2s), .qb(),
		.d(n3020), .sdi(n2212), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__23__slave ( .q(_RegFile_22__23), .qb(n2213),
		.d(_RegFile_reg_22__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__24__master ( .q(_RegFile_reg_22__24__m2s), .qb(),
		.d(n3021), .sdi(n2213), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__24__slave ( .q(_RegFile_22__24), .qb(n2214),
		.d(_RegFile_reg_22__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__25__master ( .q(_RegFile_reg_22__25__m2s), .qb(),
		.d(n3022), .sdi(n2214), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__25__slave ( .q(_RegFile_22__25), .qb(n2215),
		.d(_RegFile_reg_22__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__26__master ( .q(_RegFile_reg_22__26__m2s), .qb(),
		.d(n3023), .sdi(n2215), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__26__slave ( .q(_RegFile_22__26), .qb(n2216),
		.d(_RegFile_reg_22__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__27__master ( .q(_RegFile_reg_22__27__m2s), .qb(),
		.d(n3024), .sdi(n2216), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__27__slave ( .q(_RegFile_22__27), .qb(n2217),
		.d(_RegFile_reg_22__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__28__master ( .q(_RegFile_reg_22__28__m2s), .qb(),
		.d(n3025), .sdi(n2217), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__28__slave ( .q(_RegFile_22__28), .qb(n2218),
		.d(_RegFile_reg_22__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__29__master ( .q(_RegFile_reg_22__29__m2s), .qb(),
		.d(n3026), .sdi(n2218), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__29__slave ( .q(_RegFile_22__29), .qb(n2219),
		.d(_RegFile_reg_22__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__2__master ( .q(_RegFile_reg_22__2__m2s), .qb(),
		.d(n2999), .sdi(n4191), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__2__slave ( .q(_RegFile_22__2), .qb(n4190), .d(_RegFile_reg_22__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__30__master ( .q(_RegFile_reg_22__30__m2s), .qb(),
		.d(n3027), .sdi(n2219), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__30__slave ( .q(_RegFile_22__30), .qb(n2220),
		.d(_RegFile_reg_22__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__31__master ( .q(_RegFile_reg_22__31__m2s), .qb(),
		.d(n3028), .sdi(n2220), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__31__slave ( .q(_RegFile_22__31), .qb(n2221),
		.d(_RegFile_reg_22__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__3__master ( .q(_RegFile_reg_22__3__m2s), .qb(),
		.d(n3000), .sdi(n4190), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n936),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__3__slave ( .q(_RegFile_22__3), .qb(n4189), .d(_RegFile_reg_22__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n936), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__4__master ( .q(_RegFile_reg_22__4__m2s), .qb(),
		.d(n3001), .sdi(n4189), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__4__slave ( .q(_RegFile_22__4), .qb(n4188), .d(_RegFile_reg_22__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__5__master ( .q(_RegFile_reg_22__5__m2s), .qb(),
		.d(n3002), .sdi(n4188), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__5__slave ( .q(_RegFile_22__5), .qb(n4187), .d(_RegFile_reg_22__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__6__master ( .q(_RegFile_reg_22__6__m2s), .qb(),
		.d(n3003), .sdi(n4187), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__6__slave ( .q(_RegFile_22__6), .qb(n4186), .d(_RegFile_reg_22__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__7__master ( .q(_RegFile_reg_22__7__m2s), .qb(),
		.d(n3004), .sdi(n4186), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__7__slave ( .q(_RegFile_22__7), .qb(n4185), .d(_RegFile_reg_22__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__8__master ( .q(_RegFile_reg_22__8__m2s), .qb(),
		.d(n3005), .sdi(n4185), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__8__slave ( .q(_RegFile_22__8), .qb(n2222), .d(_RegFile_reg_22__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_22__9__master ( .q(_RegFile_reg_22__9__m2s), .qb(),
		.d(n3006), .sdi(n2222), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_22__9__slave ( .q(_RegFile_22__9), .qb(n2223), .d(_RegFile_reg_22__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__0__master ( .q(_RegFile_reg_23__0__m2s), .qb(),
		.d(n2965), .sdi(n2221), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__0__slave ( .q(_RegFile_23__0), .qb(n4184), .d(_RegFile_reg_23__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__10__master ( .q(_RegFile_reg_23__10__m2s), .qb(),
		.d(n2975), .sdi(n2247), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__10__slave ( .q(_RegFile_23__10), .qb(n2224),
		.d(_RegFile_reg_23__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__11__master ( .q(_RegFile_reg_23__11__m2s), .qb(),
		.d(n2976), .sdi(n2224), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__11__slave ( .q(_RegFile_23__11), .qb(n2225),
		.d(_RegFile_reg_23__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__12__master ( .q(_RegFile_reg_23__12__m2s), .qb(),
		.d(n2977), .sdi(n2225), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__12__slave ( .q(_RegFile_23__12), .qb(n2226),
		.d(_RegFile_reg_23__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__13__master ( .q(_RegFile_reg_23__13__m2s), .qb(),
		.d(n2978), .sdi(n2226), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__13__slave ( .q(_RegFile_23__13), .qb(n2227),
		.d(_RegFile_reg_23__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__14__master ( .q(_RegFile_reg_23__14__m2s), .qb(),
		.d(n2979), .sdi(n2227), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n966),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__14__slave ( .q(_RegFile_23__14), .qb(n2228),
		.d(_RegFile_reg_23__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n966), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__15__master ( .q(_RegFile_reg_23__15__m2s), .qb(),
		.d(n2980), .sdi(n2228), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__15__slave ( .q(_RegFile_23__15), .qb(n2229),
		.d(_RegFile_reg_23__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__16__master ( .q(_RegFile_reg_23__16__m2s), .qb(),
		.d(n2981), .sdi(n2229), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__16__slave ( .q(_RegFile_23__16), .qb(n2230),
		.d(_RegFile_reg_23__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__17__master ( .q(_RegFile_reg_23__17__m2s), .qb(),
		.d(n2982), .sdi(n2230), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__17__slave ( .q(_RegFile_23__17), .qb(n2231),
		.d(_RegFile_reg_23__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__18__master ( .q(_RegFile_reg_23__18__m2s), .qb(),
		.d(n2983), .sdi(n2231), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__18__slave ( .q(_RegFile_23__18), .qb(n2232),
		.d(_RegFile_reg_23__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__19__master ( .q(_RegFile_reg_23__19__m2s), .qb(),
		.d(n2984), .sdi(n2232), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__19__slave ( .q(_RegFile_23__19), .qb(n2233),
		.d(_RegFile_reg_23__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__1__master ( .q(_RegFile_reg_23__1__m2s), .qb(),
		.d(n2966), .sdi(n4184), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__1__slave ( .q(_RegFile_23__1), .qb(n4183), .d(_RegFile_reg_23__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__20__master ( .q(_RegFile_reg_23__20__m2s), .qb(),
		.d(n2985), .sdi(n2233), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__20__slave ( .q(_RegFile_23__20), .qb(n2234),
		.d(_RegFile_reg_23__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__21__master ( .q(_RegFile_reg_23__21__m2s), .qb(),
		.d(n2986), .sdi(n2234), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__21__slave ( .q(_RegFile_23__21), .qb(n2235),
		.d(_RegFile_reg_23__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__22__master ( .q(_RegFile_reg_23__22__m2s), .qb(),
		.d(n2987), .sdi(n2235), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__22__slave ( .q(_RegFile_23__22), .qb(n2236),
		.d(_RegFile_reg_23__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__23__master ( .q(_RegFile_reg_23__23__m2s), .qb(),
		.d(n2988), .sdi(n2236), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__23__slave ( .q(_RegFile_23__23), .qb(n2237),
		.d(_RegFile_reg_23__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__24__master ( .q(_RegFile_reg_23__24__m2s), .qb(),
		.d(n2989), .sdi(n2237), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__24__slave ( .q(_RegFile_23__24), .qb(n2238),
		.d(_RegFile_reg_23__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__25__master ( .q(_RegFile_reg_23__25__m2s), .qb(),
		.d(n2990), .sdi(n2238), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__25__slave ( .q(_RegFile_23__25), .qb(n2239),
		.d(_RegFile_reg_23__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__26__master ( .q(_RegFile_reg_23__26__m2s), .qb(),
		.d(n2991), .sdi(n2239), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__26__slave ( .q(_RegFile_23__26), .qb(n2240),
		.d(_RegFile_reg_23__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__27__master ( .q(_RegFile_reg_23__27__m2s), .qb(),
		.d(n2992), .sdi(n2240), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__27__slave ( .q(_RegFile_23__27), .qb(n2241),
		.d(_RegFile_reg_23__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__28__master ( .q(_RegFile_reg_23__28__m2s), .qb(),
		.d(n2993), .sdi(n2241), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__28__slave ( .q(_RegFile_23__28), .qb(n2242),
		.d(_RegFile_reg_23__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__29__master ( .q(_RegFile_reg_23__29__m2s), .qb(),
		.d(n2994), .sdi(n2242), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__29__slave ( .q(_RegFile_23__29), .qb(n2243),
		.d(_RegFile_reg_23__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__2__master ( .q(_RegFile_reg_23__2__m2s), .qb(),
		.d(n2967), .sdi(n4183), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__2__slave ( .q(_RegFile_23__2), .qb(n4182), .d(_RegFile_reg_23__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__30__master ( .q(_RegFile_reg_23__30__m2s), .qb(),
		.d(n2995), .sdi(n2243), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__30__slave ( .q(_RegFile_23__30), .qb(n2244),
		.d(_RegFile_reg_23__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__31__master ( .q(_RegFile_reg_23__31__m2s), .qb(),
		.d(n2996), .sdi(n2244), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__31__slave ( .q(_RegFile_23__31), .qb(n2245),
		.d(_RegFile_reg_23__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__3__master ( .q(_RegFile_reg_23__3__m2s), .qb(),
		.d(n2968), .sdi(n4182), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__3__slave ( .q(_RegFile_23__3), .qb(n4181), .d(_RegFile_reg_23__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__4__master ( .q(_RegFile_reg_23__4__m2s), .qb(),
		.d(n2969), .sdi(n4181), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__4__slave ( .q(_RegFile_23__4), .qb(n4180), .d(_RegFile_reg_23__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__5__master ( .q(_RegFile_reg_23__5__m2s), .qb(),
		.d(n2970), .sdi(n4180), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__5__slave ( .q(_RegFile_23__5), .qb(n4179), .d(_RegFile_reg_23__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__6__master ( .q(_RegFile_reg_23__6__m2s), .qb(),
		.d(n2971), .sdi(n4179), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__6__slave ( .q(_RegFile_23__6), .qb(n4178), .d(_RegFile_reg_23__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__7__master ( .q(_RegFile_reg_23__7__m2s), .qb(),
		.d(n2972), .sdi(n4178), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__7__slave ( .q(_RegFile_23__7), .qb(n4177), .d(_RegFile_reg_23__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__8__master ( .q(_RegFile_reg_23__8__m2s), .qb(),
		.d(n2973), .sdi(n4177), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__8__slave ( .q(_RegFile_23__8), .qb(n2246), .d(_RegFile_reg_23__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_23__9__master ( .q(_RegFile_reg_23__9__m2s), .qb(),
		.d(n2974), .sdi(n2246), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_23__9__slave ( .q(_RegFile_23__9), .qb(n2247), .d(_RegFile_reg_23__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__0__master ( .q(_RegFile_reg_24__0__m2s), .qb(),
		.d(n2933), .sdi(n2245), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__0__slave ( .q(_RegFile_24__0), .qb(n4176), .d(_RegFile_reg_24__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__10__master ( .q(_RegFile_reg_24__10__m2s), .qb(),
		.d(n2943), .sdi(n2271), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__10__slave ( .q(_RegFile_24__10), .qb(n2248),
		.d(_RegFile_reg_24__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__11__master ( .q(_RegFile_reg_24__11__m2s), .qb(),
		.d(n2944), .sdi(n2248), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__11__slave ( .q(_RegFile_24__11), .qb(n2249),
		.d(_RegFile_reg_24__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__12__master ( .q(_RegFile_reg_24__12__m2s), .qb(),
		.d(n2945), .sdi(n2249), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n967),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__12__slave ( .q(_RegFile_24__12), .qb(n2250),
		.d(_RegFile_reg_24__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n967), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__13__master ( .q(_RegFile_reg_24__13__m2s), .qb(),
		.d(n2946), .sdi(n2250), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__13__slave ( .q(_RegFile_24__13), .qb(n2251),
		.d(_RegFile_reg_24__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__14__master ( .q(_RegFile_reg_24__14__m2s), .qb(),
		.d(n2947), .sdi(n2251), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__14__slave ( .q(_RegFile_24__14), .qb(n2252),
		.d(_RegFile_reg_24__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__15__master ( .q(_RegFile_reg_24__15__m2s), .qb(),
		.d(n2948), .sdi(n2252), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__15__slave ( .q(_RegFile_24__15), .qb(n2253),
		.d(_RegFile_reg_24__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__16__master ( .q(_RegFile_reg_24__16__m2s), .qb(),
		.d(n2949), .sdi(n2253), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__16__slave ( .q(_RegFile_24__16), .qb(n2254),
		.d(_RegFile_reg_24__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__17__master ( .q(_RegFile_reg_24__17__m2s), .qb(),
		.d(n2950), .sdi(n2254), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__17__slave ( .q(_RegFile_24__17), .qb(n2255),
		.d(_RegFile_reg_24__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__18__master ( .q(_RegFile_reg_24__18__m2s), .qb(),
		.d(n2951), .sdi(n2255), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__18__slave ( .q(_RegFile_24__18), .qb(n2256),
		.d(_RegFile_reg_24__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__19__master ( .q(_RegFile_reg_24__19__m2s), .qb(),
		.d(n2952), .sdi(n2256), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__19__slave ( .q(_RegFile_24__19), .qb(n2257),
		.d(_RegFile_reg_24__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__1__master ( .q(_RegFile_reg_24__1__m2s), .qb(),
		.d(n2934), .sdi(n4176), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__1__slave ( .q(_RegFile_24__1), .qb(n4175), .d(_RegFile_reg_24__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__20__master ( .q(_RegFile_reg_24__20__m2s), .qb(),
		.d(n2953), .sdi(n2257), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__20__slave ( .q(_RegFile_24__20), .qb(n2258),
		.d(_RegFile_reg_24__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__21__master ( .q(_RegFile_reg_24__21__m2s), .qb(),
		.d(n2954), .sdi(n2258), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__21__slave ( .q(_RegFile_24__21), .qb(n2259),
		.d(_RegFile_reg_24__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__22__master ( .q(_RegFile_reg_24__22__m2s), .qb(),
		.d(n2955), .sdi(n2259), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__22__slave ( .q(_RegFile_24__22), .qb(n2260),
		.d(_RegFile_reg_24__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__23__master ( .q(_RegFile_reg_24__23__m2s), .qb(),
		.d(n2956), .sdi(n2260), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__23__slave ( .q(_RegFile_24__23), .qb(n2261),
		.d(_RegFile_reg_24__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__24__master ( .q(_RegFile_reg_24__24__m2s), .qb(),
		.d(n2957), .sdi(n2261), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__24__slave ( .q(_RegFile_24__24), .qb(n2262),
		.d(_RegFile_reg_24__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__25__master ( .q(_RegFile_reg_24__25__m2s), .qb(),
		.d(n2958), .sdi(n2262), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__25__slave ( .q(_RegFile_24__25), .qb(n2263),
		.d(_RegFile_reg_24__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__26__master ( .q(_RegFile_reg_24__26__m2s), .qb(),
		.d(n2959), .sdi(n2263), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n935),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__26__slave ( .q(_RegFile_24__26), .qb(n2264),
		.d(_RegFile_reg_24__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n935), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__27__master ( .q(_RegFile_reg_24__27__m2s), .qb(),
		.d(n2960), .sdi(n2264), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__27__slave ( .q(_RegFile_24__27), .qb(n2265),
		.d(_RegFile_reg_24__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__28__master ( .q(_RegFile_reg_24__28__m2s), .qb(),
		.d(n2961), .sdi(n2265), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__28__slave ( .q(_RegFile_24__28), .qb(n2266),
		.d(_RegFile_reg_24__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__29__master ( .q(_RegFile_reg_24__29__m2s), .qb(),
		.d(n2962), .sdi(n2266), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__29__slave ( .q(_RegFile_24__29), .qb(n2267),
		.d(_RegFile_reg_24__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__2__master ( .q(_RegFile_reg_24__2__m2s), .qb(),
		.d(n2935), .sdi(n4175), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__2__slave ( .q(_RegFile_24__2), .qb(n4174), .d(_RegFile_reg_24__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__30__master ( .q(_RegFile_reg_24__30__m2s), .qb(),
		.d(n2963), .sdi(n2267), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__30__slave ( .q(_RegFile_24__30), .qb(n2268),
		.d(_RegFile_reg_24__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__31__master ( .q(_RegFile_reg_24__31__m2s), .qb(),
		.d(n2964), .sdi(n2268), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__31__slave ( .q(_RegFile_24__31), .qb(n2269),
		.d(_RegFile_reg_24__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__3__master ( .q(_RegFile_reg_24__3__m2s), .qb(),
		.d(n2936), .sdi(n4174), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__3__slave ( .q(_RegFile_24__3), .qb(n4173), .d(_RegFile_reg_24__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__4__master ( .q(_RegFile_reg_24__4__m2s), .qb(),
		.d(n2937), .sdi(n4173), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__4__slave ( .q(_RegFile_24__4), .qb(n4172), .d(_RegFile_reg_24__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__5__master ( .q(_RegFile_reg_24__5__m2s), .qb(),
		.d(n2938), .sdi(n4172), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__5__slave ( .q(_RegFile_24__5), .qb(n4171), .d(_RegFile_reg_24__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__6__master ( .q(_RegFile_reg_24__6__m2s), .qb(),
		.d(n2939), .sdi(n4171), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__6__slave ( .q(_RegFile_24__6), .qb(n4170), .d(_RegFile_reg_24__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__7__master ( .q(_RegFile_reg_24__7__m2s), .qb(),
		.d(n2940), .sdi(n4170), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__7__slave ( .q(_RegFile_24__7), .qb(n4169), .d(_RegFile_reg_24__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__8__master ( .q(_RegFile_reg_24__8__m2s), .qb(),
		.d(n2941), .sdi(n4169), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__8__slave ( .q(_RegFile_24__8), .qb(n2270), .d(_RegFile_reg_24__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_24__9__master ( .q(_RegFile_reg_24__9__m2s), .qb(),
		.d(n2942), .sdi(n2270), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_24__9__slave ( .q(_RegFile_24__9), .qb(n2271), .d(_RegFile_reg_24__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__0__master ( .q(_RegFile_reg_25__0__m2s), .qb(),
		.d(n2901), .sdi(n2269), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__0__slave ( .q(_RegFile_25__0), .qb(n4168), .d(_RegFile_reg_25__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__10__master ( .q(_RegFile_reg_25__10__m2s), .qb(),
		.d(n2911), .sdi(n2295), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__10__slave ( .q(_RegFile_25__10), .qb(n2272),
		.d(_RegFile_reg_25__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__11__master ( .q(_RegFile_reg_25__11__m2s), .qb(),
		.d(n2912), .sdi(n2272), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__11__slave ( .q(_RegFile_25__11), .qb(n2273),
		.d(_RegFile_reg_25__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__12__master ( .q(_RegFile_reg_25__12__m2s), .qb(),
		.d(n2913), .sdi(n2273), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__12__slave ( .q(_RegFile_25__12), .qb(n2274),
		.d(_RegFile_reg_25__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__13__master ( .q(_RegFile_reg_25__13__m2s), .qb(),
		.d(n2914), .sdi(n2274), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__13__slave ( .q(_RegFile_25__13), .qb(n2275),
		.d(_RegFile_reg_25__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__14__master ( .q(_RegFile_reg_25__14__m2s), .qb(),
		.d(n2915), .sdi(n2275), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__14__slave ( .q(_RegFile_25__14), .qb(n2276),
		.d(_RegFile_reg_25__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__15__master ( .q(_RegFile_reg_25__15__m2s), .qb(),
		.d(n2916), .sdi(n2276), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__15__slave ( .q(_RegFile_25__15), .qb(n2277),
		.d(_RegFile_reg_25__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__16__master ( .q(_RegFile_reg_25__16__m2s), .qb(),
		.d(n2917), .sdi(n2277), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__16__slave ( .q(_RegFile_25__16), .qb(n2278),
		.d(_RegFile_reg_25__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__17__master ( .q(_RegFile_reg_25__17__m2s), .qb(),
		.d(n2918), .sdi(n2278), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__17__slave ( .q(_RegFile_25__17), .qb(n2279),
		.d(_RegFile_reg_25__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__18__master ( .q(_RegFile_reg_25__18__m2s), .qb(),
		.d(n2919), .sdi(n2279), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__18__slave ( .q(_RegFile_25__18), .qb(n2280),
		.d(_RegFile_reg_25__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__19__master ( .q(_RegFile_reg_25__19__m2s), .qb(),
		.d(n2920), .sdi(n2280), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__19__slave ( .q(_RegFile_25__19), .qb(n2281),
		.d(_RegFile_reg_25__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__1__master ( .q(_RegFile_reg_25__1__m2s), .qb(),
		.d(n2902), .sdi(n4168), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__1__slave ( .q(_RegFile_25__1), .qb(n4167), .d(_RegFile_reg_25__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__20__master ( .q(_RegFile_reg_25__20__m2s), .qb(),
		.d(n2921), .sdi(n2281), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__20__slave ( .q(_RegFile_25__20), .qb(n2282),
		.d(_RegFile_reg_25__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__21__master ( .q(_RegFile_reg_25__21__m2s), .qb(),
		.d(n2922), .sdi(n2282), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__21__slave ( .q(_RegFile_25__21), .qb(n2283),
		.d(_RegFile_reg_25__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__22__master ( .q(_RegFile_reg_25__22__m2s), .qb(),
		.d(n2923), .sdi(n2283), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__22__slave ( .q(_RegFile_25__22), .qb(n2284),
		.d(_RegFile_reg_25__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__23__master ( .q(_RegFile_reg_25__23__m2s), .qb(),
		.d(n2924), .sdi(n2284), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__23__slave ( .q(_RegFile_25__23), .qb(n2285),
		.d(_RegFile_reg_25__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__24__master ( .q(_RegFile_reg_25__24__m2s), .qb(),
		.d(n2925), .sdi(n2285), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n950),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__24__slave ( .q(_RegFile_25__24), .qb(n2286),
		.d(_RegFile_reg_25__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n950), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__25__master ( .q(_RegFile_reg_25__25__m2s), .qb(),
		.d(n2926), .sdi(n2286), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__25__slave ( .q(_RegFile_25__25), .qb(n2287),
		.d(_RegFile_reg_25__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__26__master ( .q(_RegFile_reg_25__26__m2s), .qb(),
		.d(n2927), .sdi(n2287), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__26__slave ( .q(_RegFile_25__26), .qb(n2288),
		.d(_RegFile_reg_25__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__27__master ( .q(_RegFile_reg_25__27__m2s), .qb(),
		.d(n2928), .sdi(n2288), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__27__slave ( .q(_RegFile_25__27), .qb(n2289),
		.d(_RegFile_reg_25__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__28__master ( .q(_RegFile_reg_25__28__m2s), .qb(),
		.d(n2929), .sdi(n2289), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__28__slave ( .q(_RegFile_25__28), .qb(n2290),
		.d(_RegFile_reg_25__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__29__master ( .q(_RegFile_reg_25__29__m2s), .qb(),
		.d(n2930), .sdi(n2290), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__29__slave ( .q(_RegFile_25__29), .qb(n2291),
		.d(_RegFile_reg_25__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__2__master ( .q(_RegFile_reg_25__2__m2s), .qb(),
		.d(n2903), .sdi(n4167), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__2__slave ( .q(_RegFile_25__2), .qb(n4166), .d(_RegFile_reg_25__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__30__master ( .q(_RegFile_reg_25__30__m2s), .qb(),
		.d(n2931), .sdi(n2291), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__30__slave ( .q(_RegFile_25__30), .qb(n2292),
		.d(_RegFile_reg_25__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__31__master ( .q(_RegFile_reg_25__31__m2s), .qb(),
		.d(n2932), .sdi(n2292), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__31__slave ( .q(_RegFile_25__31), .qb(n2293),
		.d(_RegFile_reg_25__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__3__master ( .q(_RegFile_reg_25__3__m2s), .qb(),
		.d(n2904), .sdi(n4166), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__3__slave ( .q(_RegFile_25__3), .qb(n4165), .d(_RegFile_reg_25__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__4__master ( .q(_RegFile_reg_25__4__m2s), .qb(),
		.d(n2905), .sdi(n4165), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__4__slave ( .q(_RegFile_25__4), .qb(n4164), .d(_RegFile_reg_25__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__5__master ( .q(_RegFile_reg_25__5__m2s), .qb(),
		.d(n2906), .sdi(n4164), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__5__slave ( .q(_RegFile_25__5), .qb(n4163), .d(_RegFile_reg_25__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__6__master ( .q(_RegFile_reg_25__6__m2s), .qb(),
		.d(n2907), .sdi(n4163), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__6__slave ( .q(_RegFile_25__6), .qb(n4162), .d(_RegFile_reg_25__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__7__master ( .q(_RegFile_reg_25__7__m2s), .qb(),
		.d(n2908), .sdi(n4162), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__7__slave ( .q(_RegFile_25__7), .qb(n4161), .d(_RegFile_reg_25__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__8__master ( .q(_RegFile_reg_25__8__m2s), .qb(),
		.d(n2909), .sdi(n4161), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__8__slave ( .q(_RegFile_25__8), .qb(n2294), .d(_RegFile_reg_25__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_25__9__master ( .q(_RegFile_reg_25__9__m2s), .qb(),
		.d(n2910), .sdi(n2294), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_25__9__slave ( .q(_RegFile_25__9), .qb(n2295), .d(_RegFile_reg_25__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__0__master ( .q(_RegFile_reg_26__0__m2s), .qb(),
		.d(n2869), .sdi(n2293), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__0__slave ( .q(_RegFile_26__0), .qb(n4160), .d(_RegFile_reg_26__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__10__master ( .q(_RegFile_reg_26__10__m2s), .qb(),
		.d(n2879), .sdi(n2319), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__10__slave ( .q(_RegFile_26__10), .qb(n2296),
		.d(_RegFile_reg_26__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__11__master ( .q(_RegFile_reg_26__11__m2s), .qb(),
		.d(n2880), .sdi(n2296), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__11__slave ( .q(_RegFile_26__11), .qb(n2297),
		.d(_RegFile_reg_26__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__12__master ( .q(_RegFile_reg_26__12__m2s), .qb(),
		.d(n2881), .sdi(n2297), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__12__slave ( .q(_RegFile_26__12), .qb(n2298),
		.d(_RegFile_reg_26__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__13__master ( .q(_RegFile_reg_26__13__m2s), .qb(),
		.d(n2882), .sdi(n2298), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__13__slave ( .q(_RegFile_26__13), .qb(n2299),
		.d(_RegFile_reg_26__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__14__master ( .q(_RegFile_reg_26__14__m2s), .qb(),
		.d(n2883), .sdi(n2299), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__14__slave ( .q(_RegFile_26__14), .qb(n2300),
		.d(_RegFile_reg_26__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__15__master ( .q(_RegFile_reg_26__15__m2s), .qb(),
		.d(n2884), .sdi(n2300), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__15__slave ( .q(_RegFile_26__15), .qb(n2301),
		.d(_RegFile_reg_26__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__16__master ( .q(_RegFile_reg_26__16__m2s), .qb(),
		.d(n2885), .sdi(n2301), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__16__slave ( .q(_RegFile_26__16), .qb(n2302),
		.d(_RegFile_reg_26__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__17__master ( .q(_RegFile_reg_26__17__m2s), .qb(),
		.d(n2886), .sdi(n2302), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__17__slave ( .q(_RegFile_26__17), .qb(n2303),
		.d(_RegFile_reg_26__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__18__master ( .q(_RegFile_reg_26__18__m2s), .qb(),
		.d(n2887), .sdi(n2303), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__18__slave ( .q(_RegFile_26__18), .qb(n2304),
		.d(_RegFile_reg_26__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__19__master ( .q(_RegFile_reg_26__19__m2s), .qb(),
		.d(n2888), .sdi(n2304), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__19__slave ( .q(_RegFile_26__19), .qb(n2305),
		.d(_RegFile_reg_26__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__1__master ( .q(_RegFile_reg_26__1__m2s), .qb(),
		.d(n2870), .sdi(n4160), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__1__slave ( .q(_RegFile_26__1), .qb(n4159), .d(_RegFile_reg_26__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__20__master ( .q(_RegFile_reg_26__20__m2s), .qb(),
		.d(n2889), .sdi(n2305), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__20__slave ( .q(_RegFile_26__20), .qb(n2306),
		.d(_RegFile_reg_26__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__21__master ( .q(_RegFile_reg_26__21__m2s), .qb(),
		.d(n2890), .sdi(n2306), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__21__slave ( .q(_RegFile_26__21), .qb(n2307),
		.d(_RegFile_reg_26__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__22__master ( .q(_RegFile_reg_26__22__m2s), .qb(),
		.d(n2891), .sdi(n2307), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n934),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__22__slave ( .q(_RegFile_26__22), .qb(n2308),
		.d(_RegFile_reg_26__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n934), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__23__master ( .q(_RegFile_reg_26__23__m2s), .qb(),
		.d(n2892), .sdi(n2308), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__23__slave ( .q(_RegFile_26__23), .qb(n2309),
		.d(_RegFile_reg_26__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__24__master ( .q(_RegFile_reg_26__24__m2s), .qb(),
		.d(n2893), .sdi(n2309), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__24__slave ( .q(_RegFile_26__24), .qb(n2310),
		.d(_RegFile_reg_26__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__25__master ( .q(_RegFile_reg_26__25__m2s), .qb(),
		.d(n2894), .sdi(n2310), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__25__slave ( .q(_RegFile_26__25), .qb(n2311),
		.d(_RegFile_reg_26__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__26__master ( .q(_RegFile_reg_26__26__m2s), .qb(),
		.d(n2895), .sdi(n2311), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__26__slave ( .q(_RegFile_26__26), .qb(n2312),
		.d(_RegFile_reg_26__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__27__master ( .q(_RegFile_reg_26__27__m2s), .qb(),
		.d(n2896), .sdi(n2312), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__27__slave ( .q(_RegFile_26__27), .qb(n2313),
		.d(_RegFile_reg_26__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__28__master ( .q(_RegFile_reg_26__28__m2s), .qb(),
		.d(n2897), .sdi(n2313), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__28__slave ( .q(_RegFile_26__28), .qb(n2314),
		.d(_RegFile_reg_26__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__29__master ( .q(_RegFile_reg_26__29__m2s), .qb(),
		.d(n2898), .sdi(n2314), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__29__slave ( .q(_RegFile_26__29), .qb(n2315),
		.d(_RegFile_reg_26__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__2__master ( .q(_RegFile_reg_26__2__m2s), .qb(),
		.d(n2871), .sdi(n4159), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__2__slave ( .q(_RegFile_26__2), .qb(n4158), .d(_RegFile_reg_26__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__30__master ( .q(_RegFile_reg_26__30__m2s), .qb(),
		.d(n2899), .sdi(n2315), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__30__slave ( .q(_RegFile_26__30), .qb(n2316),
		.d(_RegFile_reg_26__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__31__master ( .q(_RegFile_reg_26__31__m2s), .qb(),
		.d(n2900), .sdi(n2316), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__31__slave ( .q(_RegFile_26__31), .qb(n2317),
		.d(_RegFile_reg_26__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__3__master ( .q(_RegFile_reg_26__3__m2s), .qb(),
		.d(n2872), .sdi(n4158), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__3__slave ( .q(_RegFile_26__3), .qb(n4157), .d(_RegFile_reg_26__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__4__master ( .q(_RegFile_reg_26__4__m2s), .qb(),
		.d(n2873), .sdi(n4157), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__4__slave ( .q(_RegFile_26__4), .qb(n4156), .d(_RegFile_reg_26__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__5__master ( .q(_RegFile_reg_26__5__m2s), .qb(),
		.d(n2874), .sdi(n4156), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__5__slave ( .q(_RegFile_26__5), .qb(n4155), .d(_RegFile_reg_26__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__6__master ( .q(_RegFile_reg_26__6__m2s), .qb(),
		.d(n2875), .sdi(n4155), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__6__slave ( .q(_RegFile_26__6), .qb(n4154), .d(_RegFile_reg_26__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__7__master ( .q(_RegFile_reg_26__7__m2s), .qb(),
		.d(n2876), .sdi(n4154), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__7__slave ( .q(_RegFile_26__7), .qb(n4153), .d(_RegFile_reg_26__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__8__master ( .q(_RegFile_reg_26__8__m2s), .qb(),
		.d(n2877), .sdi(n4153), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n970),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__8__slave ( .q(_RegFile_26__8), .qb(n2318), .d(_RegFile_reg_26__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n970), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_26__9__master ( .q(_RegFile_reg_26__9__m2s), .qb(),
		.d(n2878), .sdi(n2318), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_26__9__slave ( .q(_RegFile_26__9), .qb(n2319), .d(_RegFile_reg_26__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__0__master ( .q(_RegFile_reg_27__0__m2s), .qb(),
		.d(n2837), .sdi(n2317), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__0__slave ( .q(_RegFile_27__0), .qb(n4152), .d(_RegFile_reg_27__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__10__master ( .q(_RegFile_reg_27__10__m2s), .qb(),
		.d(n2847), .sdi(n2343), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__10__slave ( .q(_RegFile_27__10), .qb(n2320),
		.d(_RegFile_reg_27__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__11__master ( .q(_RegFile_reg_27__11__m2s), .qb(),
		.d(n2848), .sdi(n2320), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__11__slave ( .q(_RegFile_27__11), .qb(n2321),
		.d(_RegFile_reg_27__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__12__master ( .q(_RegFile_reg_27__12__m2s), .qb(),
		.d(n2849), .sdi(n2321), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__12__slave ( .q(_RegFile_27__12), .qb(n2322),
		.d(_RegFile_reg_27__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__13__master ( .q(_RegFile_reg_27__13__m2s), .qb(),
		.d(n2850), .sdi(n2322), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__13__slave ( .q(_RegFile_27__13), .qb(n2323),
		.d(_RegFile_reg_27__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__14__master ( .q(_RegFile_reg_27__14__m2s), .qb(),
		.d(n2851), .sdi(n2323), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__14__slave ( .q(_RegFile_27__14), .qb(n2324),
		.d(_RegFile_reg_27__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__15__master ( .q(_RegFile_reg_27__15__m2s), .qb(),
		.d(n2852), .sdi(n2324), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__15__slave ( .q(_RegFile_27__15), .qb(n2325),
		.d(_RegFile_reg_27__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__16__master ( .q(_RegFile_reg_27__16__m2s), .qb(),
		.d(n2853), .sdi(n2325), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__16__slave ( .q(_RegFile_27__16), .qb(n2326),
		.d(_RegFile_reg_27__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__17__master ( .q(_RegFile_reg_27__17__m2s), .qb(),
		.d(n2854), .sdi(n2326), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__17__slave ( .q(_RegFile_27__17), .qb(n2327),
		.d(_RegFile_reg_27__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__18__master ( .q(_RegFile_reg_27__18__m2s), .qb(),
		.d(n2855), .sdi(n2327), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__18__slave ( .q(_RegFile_27__18), .qb(n2328),
		.d(_RegFile_reg_27__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__19__master ( .q(_RegFile_reg_27__19__m2s), .qb(),
		.d(n2856), .sdi(n2328), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__19__slave ( .q(_RegFile_27__19), .qb(n2329),
		.d(_RegFile_reg_27__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__1__master ( .q(_RegFile_reg_27__1__m2s), .qb(),
		.d(n2838), .sdi(n4152), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__1__slave ( .q(_RegFile_27__1), .qb(n4151), .d(_RegFile_reg_27__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__20__master ( .q(_RegFile_reg_27__20__m2s), .qb(),
		.d(n2857), .sdi(n2329), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n933),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__20__slave ( .q(_RegFile_27__20), .qb(n2330),
		.d(_RegFile_reg_27__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n933), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__21__master ( .q(_RegFile_reg_27__21__m2s), .qb(),
		.d(n2858), .sdi(n2330), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__21__slave ( .q(_RegFile_27__21), .qb(n2331),
		.d(_RegFile_reg_27__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__22__master ( .q(_RegFile_reg_27__22__m2s), .qb(),
		.d(n2859), .sdi(n2331), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__22__slave ( .q(_RegFile_27__22), .qb(n2332),
		.d(_RegFile_reg_27__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__23__master ( .q(_RegFile_reg_27__23__m2s), .qb(),
		.d(n2860), .sdi(n2332), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__23__slave ( .q(_RegFile_27__23), .qb(n2333),
		.d(_RegFile_reg_27__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__24__master ( .q(_RegFile_reg_27__24__m2s), .qb(),
		.d(n2861), .sdi(n2333), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__24__slave ( .q(_RegFile_27__24), .qb(n2334),
		.d(_RegFile_reg_27__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__25__master ( .q(_RegFile_reg_27__25__m2s), .qb(),
		.d(n2862), .sdi(n2334), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__25__slave ( .q(_RegFile_27__25), .qb(n2335),
		.d(_RegFile_reg_27__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__26__master ( .q(_RegFile_reg_27__26__m2s), .qb(),
		.d(n2863), .sdi(n2335), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__26__slave ( .q(_RegFile_27__26), .qb(n2336),
		.d(_RegFile_reg_27__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__27__master ( .q(_RegFile_reg_27__27__m2s), .qb(),
		.d(n2864), .sdi(n2336), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__27__slave ( .q(_RegFile_27__27), .qb(n2337),
		.d(_RegFile_reg_27__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__28__master ( .q(_RegFile_reg_27__28__m2s), .qb(),
		.d(n2865), .sdi(n2337), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__28__slave ( .q(_RegFile_27__28), .qb(n2338),
		.d(_RegFile_reg_27__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__29__master ( .q(_RegFile_reg_27__29__m2s), .qb(),
		.d(n2866), .sdi(n2338), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__29__slave ( .q(_RegFile_27__29), .qb(n2339),
		.d(_RegFile_reg_27__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__2__master ( .q(_RegFile_reg_27__2__m2s), .qb(),
		.d(n2839), .sdi(n4151), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__2__slave ( .q(_RegFile_27__2), .qb(n4150), .d(_RegFile_reg_27__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__30__master ( .q(_RegFile_reg_27__30__m2s), .qb(),
		.d(n2867), .sdi(n2339), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__30__slave ( .q(_RegFile_27__30), .qb(n2340),
		.d(_RegFile_reg_27__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__31__master ( .q(_RegFile_reg_27__31__m2s), .qb(),
		.d(n2868), .sdi(n2340), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__31__slave ( .q(_RegFile_27__31), .qb(n2341),
		.d(_RegFile_reg_27__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__3__master ( .q(_RegFile_reg_27__3__m2s), .qb(),
		.d(n2840), .sdi(n4150), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__3__slave ( .q(_RegFile_27__3), .qb(n4149), .d(_RegFile_reg_27__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__4__master ( .q(_RegFile_reg_27__4__m2s), .qb(),
		.d(n2841), .sdi(n4149), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__4__slave ( .q(_RegFile_27__4), .qb(n4148), .d(_RegFile_reg_27__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__5__master ( .q(_RegFile_reg_27__5__m2s), .qb(),
		.d(n2842), .sdi(n4148), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__5__slave ( .q(_RegFile_27__5), .qb(n4147), .d(_RegFile_reg_27__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__6__master ( .q(_RegFile_reg_27__6__m2s), .qb(),
		.d(n2843), .sdi(n4147), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n971),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__6__slave ( .q(_RegFile_27__6), .qb(n4146), .d(_RegFile_reg_27__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n971), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__7__master ( .q(_RegFile_reg_27__7__m2s), .qb(),
		.d(n2844), .sdi(n4146), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__7__slave ( .q(_RegFile_27__7), .qb(n4145), .d(_RegFile_reg_27__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__8__master ( .q(_RegFile_reg_27__8__m2s), .qb(),
		.d(n2845), .sdi(n4145), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__8__slave ( .q(_RegFile_27__8), .qb(n2342), .d(_RegFile_reg_27__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_27__9__master ( .q(_RegFile_reg_27__9__m2s), .qb(),
		.d(n2846), .sdi(n2342), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_27__9__slave ( .q(_RegFile_27__9), .qb(n2343), .d(_RegFile_reg_27__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__0__master ( .q(_RegFile_reg_28__0__m2s), .qb(),
		.d(n2805), .sdi(n2341), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__0__slave ( .q(_RegFile_28__0), .qb(n4144), .d(_RegFile_reg_28__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__10__master ( .q(_RegFile_reg_28__10__m2s), .qb(),
		.d(n2815), .sdi(n2367), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__10__slave ( .q(_RegFile_28__10), .qb(n2344),
		.d(_RegFile_reg_28__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__11__master ( .q(_RegFile_reg_28__11__m2s), .qb(),
		.d(n2816), .sdi(n2344), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__11__slave ( .q(_RegFile_28__11), .qb(n2345),
		.d(_RegFile_reg_28__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__12__master ( .q(_RegFile_reg_28__12__m2s), .qb(),
		.d(n2817), .sdi(n2345), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__12__slave ( .q(_RegFile_28__12), .qb(n2346),
		.d(_RegFile_reg_28__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__13__master ( .q(_RegFile_reg_28__13__m2s), .qb(),
		.d(n2818), .sdi(n2346), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__13__slave ( .q(_RegFile_28__13), .qb(n2347),
		.d(_RegFile_reg_28__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__14__master ( .q(_RegFile_reg_28__14__m2s), .qb(),
		.d(n2819), .sdi(n2347), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__14__slave ( .q(_RegFile_28__14), .qb(n2348),
		.d(_RegFile_reg_28__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__15__master ( .q(_RegFile_reg_28__15__m2s), .qb(),
		.d(n2820), .sdi(n2348), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__15__slave ( .q(_RegFile_28__15), .qb(n2349),
		.d(_RegFile_reg_28__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__16__master ( .q(_RegFile_reg_28__16__m2s), .qb(),
		.d(n2821), .sdi(n2349), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__16__slave ( .q(_RegFile_28__16), .qb(n2350),
		.d(_RegFile_reg_28__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__17__master ( .q(_RegFile_reg_28__17__m2s), .qb(),
		.d(n2822), .sdi(n2350), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__17__slave ( .q(_RegFile_28__17), .qb(n2351),
		.d(_RegFile_reg_28__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__18__master ( .q(_RegFile_reg_28__18__m2s), .qb(),
		.d(n2823), .sdi(n2351), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__18__slave ( .q(_RegFile_28__18), .qb(n2352),
		.d(_RegFile_reg_28__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__19__master ( .q(_RegFile_reg_28__19__m2s), .qb(),
		.d(n2824), .sdi(n2352), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__19__slave ( .q(_RegFile_28__19), .qb(n2353),
		.d(_RegFile_reg_28__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__1__master ( .q(_RegFile_reg_28__1__m2s), .qb(),
		.d(n2806), .sdi(n4144), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n932),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__1__slave ( .q(_RegFile_28__1), .qb(n4143), .d(_RegFile_reg_28__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n932), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__20__master ( .q(_RegFile_reg_28__20__m2s), .qb(),
		.d(n2825), .sdi(n2353), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__20__slave ( .q(_RegFile_28__20), .qb(n2354),
		.d(_RegFile_reg_28__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__21__master ( .q(_RegFile_reg_28__21__m2s), .qb(),
		.d(n2826), .sdi(n2354), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__21__slave ( .q(_RegFile_28__21), .qb(n2355),
		.d(_RegFile_reg_28__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__22__master ( .q(_RegFile_reg_28__22__m2s), .qb(),
		.d(n2827), .sdi(n2355), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__22__slave ( .q(_RegFile_28__22), .qb(n2356),
		.d(_RegFile_reg_28__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__23__master ( .q(_RegFile_reg_28__23__m2s), .qb(),
		.d(n2828), .sdi(n2356), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__23__slave ( .q(_RegFile_28__23), .qb(n2357),
		.d(_RegFile_reg_28__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__24__master ( .q(_RegFile_reg_28__24__m2s), .qb(),
		.d(n2829), .sdi(n2357), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__24__slave ( .q(_RegFile_28__24), .qb(n2358),
		.d(_RegFile_reg_28__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__25__master ( .q(_RegFile_reg_28__25__m2s), .qb(),
		.d(n2830), .sdi(n2358), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__25__slave ( .q(_RegFile_28__25), .qb(n2359),
		.d(_RegFile_reg_28__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__26__master ( .q(_RegFile_reg_28__26__m2s), .qb(),
		.d(n2831), .sdi(n2359), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__26__slave ( .q(_RegFile_28__26), .qb(n2360),
		.d(_RegFile_reg_28__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__27__master ( .q(_RegFile_reg_28__27__m2s), .qb(),
		.d(n2832), .sdi(n2360), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__27__slave ( .q(_RegFile_28__27), .qb(n2361),
		.d(_RegFile_reg_28__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__28__master ( .q(_RegFile_reg_28__28__m2s), .qb(),
		.d(n2833), .sdi(n2361), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__28__slave ( .q(_RegFile_28__28), .qb(n2362),
		.d(_RegFile_reg_28__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__29__master ( .q(_RegFile_reg_28__29__m2s), .qb(),
		.d(n2834), .sdi(n2362), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__29__slave ( .q(_RegFile_28__29), .qb(n2363),
		.d(_RegFile_reg_28__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__2__master ( .q(_RegFile_reg_28__2__m2s), .qb(),
		.d(n2807), .sdi(n4143), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__2__slave ( .q(_RegFile_28__2), .qb(n4142), .d(_RegFile_reg_28__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__30__master ( .q(_RegFile_reg_28__30__m2s), .qb(),
		.d(n2835), .sdi(n2363), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__30__slave ( .q(_RegFile_28__30), .qb(n2364),
		.d(_RegFile_reg_28__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__31__master ( .q(_RegFile_reg_28__31__m2s), .qb(),
		.d(n2836), .sdi(n2364), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__31__slave ( .q(_RegFile_28__31), .qb(n2365),
		.d(_RegFile_reg_28__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__3__master ( .q(_RegFile_reg_28__3__m2s), .qb(),
		.d(n2808), .sdi(n4142), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__3__slave ( .q(_RegFile_28__3), .qb(n4141), .d(_RegFile_reg_28__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__4__master ( .q(_RegFile_reg_28__4__m2s), .qb(),
		.d(n2809), .sdi(n4141), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n968),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__4__slave ( .q(_RegFile_28__4), .qb(n4140), .d(_RegFile_reg_28__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n968), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__5__master ( .q(_RegFile_reg_28__5__m2s), .qb(),
		.d(n2810), .sdi(n4140), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__5__slave ( .q(_RegFile_28__5), .qb(n4139), .d(_RegFile_reg_28__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__6__master ( .q(_RegFile_reg_28__6__m2s), .qb(),
		.d(n2811), .sdi(n4139), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__6__slave ( .q(_RegFile_28__6), .qb(n4138), .d(_RegFile_reg_28__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__7__master ( .q(_RegFile_reg_28__7__m2s), .qb(),
		.d(n2812), .sdi(n4138), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__7__slave ( .q(_RegFile_28__7), .qb(n4137), .d(_RegFile_reg_28__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__8__master ( .q(_RegFile_reg_28__8__m2s), .qb(),
		.d(n2813), .sdi(n4137), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__8__slave ( .q(_RegFile_28__8), .qb(n2366), .d(_RegFile_reg_28__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_28__9__master ( .q(_RegFile_reg_28__9__m2s), .qb(),
		.d(n2814), .sdi(n2366), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_28__9__slave ( .q(_RegFile_28__9), .qb(n2367), .d(_RegFile_reg_28__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__0__master ( .q(_RegFile_reg_29__0__m2s), .qb(),
		.d(n2773), .sdi(n2365), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__0__slave ( .q(_RegFile_29__0), .qb(n4136), .d(_RegFile_reg_29__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__10__master ( .q(_RegFile_reg_29__10__m2s), .qb(),
		.d(n2783), .sdi(n2391), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__10__slave ( .q(_RegFile_29__10), .qb(n2368),
		.d(_RegFile_reg_29__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__11__master ( .q(_RegFile_reg_29__11__m2s), .qb(),
		.d(n2784), .sdi(n2368), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__11__slave ( .q(_RegFile_29__11), .qb(n2369),
		.d(_RegFile_reg_29__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__12__master ( .q(_RegFile_reg_29__12__m2s), .qb(),
		.d(n2785), .sdi(n2369), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__12__slave ( .q(_RegFile_29__12), .qb(n2370),
		.d(_RegFile_reg_29__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__13__master ( .q(_RegFile_reg_29__13__m2s), .qb(),
		.d(n2786), .sdi(n2370), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__13__slave ( .q(_RegFile_29__13), .qb(n2371),
		.d(_RegFile_reg_29__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__14__master ( .q(_RegFile_reg_29__14__m2s), .qb(),
		.d(n2787), .sdi(n2371), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__14__slave ( .q(_RegFile_29__14), .qb(n2372),
		.d(_RegFile_reg_29__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__15__master ( .q(_RegFile_reg_29__15__m2s), .qb(),
		.d(n2788), .sdi(n2372), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__15__slave ( .q(_RegFile_29__15), .qb(n2373),
		.d(_RegFile_reg_29__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__16__master ( .q(_RegFile_reg_29__16__m2s), .qb(),
		.d(n2789), .sdi(n2373), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__16__slave ( .q(_RegFile_29__16), .qb(n2374),
		.d(_RegFile_reg_29__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__17__master ( .q(_RegFile_reg_29__17__m2s), .qb(),
		.d(n2790), .sdi(n2374), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__17__slave ( .q(_RegFile_29__17), .qb(n2375),
		.d(_RegFile_reg_29__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__18__master ( .q(_RegFile_reg_29__18__m2s), .qb(),
		.d(n2791), .sdi(n2375), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__18__slave ( .q(_RegFile_29__18), .qb(n2376),
		.d(_RegFile_reg_29__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__19__master ( .q(_RegFile_reg_29__19__m2s), .qb(),
		.d(n2792), .sdi(n2376), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__19__slave ( .q(_RegFile_29__19), .qb(n2377),
		.d(_RegFile_reg_29__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__1__master ( .q(_RegFile_reg_29__1__m2s), .qb(),
		.d(n2774), .sdi(n4136), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n931),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__1__slave ( .q(_RegFile_29__1), .qb(n4135), .d(_RegFile_reg_29__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n931), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__20__master ( .q(_RegFile_reg_29__20__m2s), .qb(),
		.d(n2793), .sdi(n2377), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__20__slave ( .q(_RegFile_29__20), .qb(n2378),
		.d(_RegFile_reg_29__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__21__master ( .q(_RegFile_reg_29__21__m2s), .qb(),
		.d(n2794), .sdi(n2378), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__21__slave ( .q(_RegFile_29__21), .qb(n2379),
		.d(_RegFile_reg_29__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__22__master ( .q(_RegFile_reg_29__22__m2s), .qb(),
		.d(n2795), .sdi(n2379), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__22__slave ( .q(_RegFile_29__22), .qb(n2380),
		.d(_RegFile_reg_29__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__23__master ( .q(_RegFile_reg_29__23__m2s), .qb(),
		.d(n2796), .sdi(n2380), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__23__slave ( .q(_RegFile_29__23), .qb(n2381),
		.d(_RegFile_reg_29__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__24__master ( .q(_RegFile_reg_29__24__m2s), .qb(),
		.d(n2797), .sdi(n2381), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__24__slave ( .q(_RegFile_29__24), .qb(n2382),
		.d(_RegFile_reg_29__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__25__master ( .q(_RegFile_reg_29__25__m2s), .qb(),
		.d(n2798), .sdi(n2382), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__25__slave ( .q(_RegFile_29__25), .qb(n2383),
		.d(_RegFile_reg_29__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__26__master ( .q(_RegFile_reg_29__26__m2s), .qb(),
		.d(n2799), .sdi(n2383), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__26__slave ( .q(_RegFile_29__26), .qb(n2384),
		.d(_RegFile_reg_29__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__27__master ( .q(_RegFile_reg_29__27__m2s), .qb(),
		.d(n2800), .sdi(n2384), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__27__slave ( .q(_RegFile_29__27), .qb(n2385),
		.d(_RegFile_reg_29__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__28__master ( .q(_RegFile_reg_29__28__m2s), .qb(),
		.d(n2801), .sdi(n2385), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__28__slave ( .q(_RegFile_29__28), .qb(n2386),
		.d(_RegFile_reg_29__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__29__master ( .q(_RegFile_reg_29__29__m2s), .qb(),
		.d(n2802), .sdi(n2386), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__29__slave ( .q(_RegFile_29__29), .qb(n2387),
		.d(_RegFile_reg_29__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__2__master ( .q(_RegFile_reg_29__2__m2s), .qb(),
		.d(n2775), .sdi(n4135), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__2__slave ( .q(_RegFile_29__2), .qb(n4134), .d(_RegFile_reg_29__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__30__master ( .q(_RegFile_reg_29__30__m2s), .qb(),
		.d(n2803), .sdi(n2387), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n972),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__30__slave ( .q(_RegFile_29__30), .qb(n2388),
		.d(_RegFile_reg_29__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n972), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__31__master ( .q(_RegFile_reg_29__31__m2s), .qb(),
		.d(n2804), .sdi(n2388), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__31__slave ( .q(_RegFile_29__31), .qb(n2389),
		.d(_RegFile_reg_29__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__3__master ( .q(_RegFile_reg_29__3__m2s), .qb(),
		.d(n2776), .sdi(n4134), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__3__slave ( .q(_RegFile_29__3), .qb(n4133), .d(_RegFile_reg_29__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__4__master ( .q(_RegFile_reg_29__4__m2s), .qb(),
		.d(n2777), .sdi(n4133), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__4__slave ( .q(_RegFile_29__4), .qb(n4132), .d(_RegFile_reg_29__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__5__master ( .q(_RegFile_reg_29__5__m2s), .qb(),
		.d(n2778), .sdi(n4132), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__5__slave ( .q(_RegFile_29__5), .qb(n4131), .d(_RegFile_reg_29__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__6__master ( .q(_RegFile_reg_29__6__m2s), .qb(),
		.d(n2779), .sdi(n4131), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__6__slave ( .q(_RegFile_29__6), .qb(n4130), .d(_RegFile_reg_29__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__7__master ( .q(_RegFile_reg_29__7__m2s), .qb(),
		.d(n2780), .sdi(n4130), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__7__slave ( .q(_RegFile_29__7), .qb(n4129), .d(_RegFile_reg_29__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__8__master ( .q(_RegFile_reg_29__8__m2s), .qb(),
		.d(n2781), .sdi(n4129), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__8__slave ( .q(_RegFile_29__8), .qb(n2390), .d(_RegFile_reg_29__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_29__9__master ( .q(_RegFile_reg_29__9__m2s), .qb(),
		.d(n2782), .sdi(n2390), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_29__9__slave ( .q(_RegFile_29__9), .qb(n2391), .d(_RegFile_reg_29__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__0__master ( .q(_RegFile_reg_2__0__m2s), .qb(),
		.d(n3637), .sdi(n2149), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__0__slave ( .q(_RegFile_2__0), .qb(n4352), .d(_RegFile_reg_2__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__10__master ( .q(_RegFile_reg_2__10__m2s), .qb(),
		.d(n3647), .sdi(n2415), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__10__slave ( .q(_RegFile_2__10), .qb(n2392), .d(_RegFile_reg_2__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__11__master ( .q(_RegFile_reg_2__11__m2s), .qb(),
		.d(n3648), .sdi(n2392), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__11__slave ( .q(_RegFile_2__11), .qb(n2393), .d(_RegFile_reg_2__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__12__master ( .q(_RegFile_reg_2__12__m2s), .qb(),
		.d(n3649), .sdi(n2393), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__12__slave ( .q(_RegFile_2__12), .qb(n2394), .d(_RegFile_reg_2__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__13__master ( .q(_RegFile_reg_2__13__m2s), .qb(),
		.d(n3650), .sdi(n2394), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__13__slave ( .q(_RegFile_2__13), .qb(n2395), .d(_RegFile_reg_2__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__14__master ( .q(_RegFile_reg_2__14__m2s), .qb(),
		.d(n3651), .sdi(n2395), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__14__slave ( .q(_RegFile_2__14), .qb(n2396), .d(_RegFile_reg_2__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__15__master ( .q(_RegFile_reg_2__15__m2s), .qb(),
		.d(n3652), .sdi(n2396), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__15__slave ( .q(_RegFile_2__15), .qb(n2397), .d(_RegFile_reg_2__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__16__master ( .q(_RegFile_reg_2__16__m2s), .qb(),
		.d(n3653), .sdi(n2397), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__16__slave ( .q(_RegFile_2__16), .qb(n2398), .d(_RegFile_reg_2__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__17__master ( .q(_RegFile_reg_2__17__m2s), .qb(),
		.d(n3654), .sdi(n2398), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__17__slave ( .q(_RegFile_2__17), .qb(n2399), .d(_RegFile_reg_2__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__18__master ( .q(_RegFile_reg_2__18__m2s), .qb(),
		.d(n3655), .sdi(n2399), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__18__slave ( .q(_RegFile_2__18), .qb(n2400), .d(_RegFile_reg_2__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__19__master ( .q(_RegFile_reg_2__19__m2s), .qb(),
		.d(n3656), .sdi(n2400), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__19__slave ( .q(_RegFile_2__19), .qb(n2401), .d(_RegFile_reg_2__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__1__master ( .q(_RegFile_reg_2__1__m2s), .qb(),
		.d(n3638), .sdi(n4352), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n930),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__1__slave ( .q(_RegFile_2__1), .qb(n4351), .d(_RegFile_reg_2__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n930), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__20__master ( .q(_RegFile_reg_2__20__m2s), .qb(),
		.d(n3657), .sdi(n2401), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__20__slave ( .q(_RegFile_2__20), .qb(n2402), .d(_RegFile_reg_2__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__21__master ( .q(_RegFile_reg_2__21__m2s), .qb(),
		.d(n3658), .sdi(n2402), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__21__slave ( .q(_RegFile_2__21), .qb(n2403), .d(_RegFile_reg_2__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__22__master ( .q(_RegFile_reg_2__22__m2s), .qb(),
		.d(n3659), .sdi(n2403), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__22__slave ( .q(_RegFile_2__22), .qb(n2404), .d(_RegFile_reg_2__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__23__master ( .q(_RegFile_reg_2__23__m2s), .qb(),
		.d(n3660), .sdi(n2404), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__23__slave ( .q(_RegFile_2__23), .qb(n2405), .d(_RegFile_reg_2__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__24__master ( .q(_RegFile_reg_2__24__m2s), .qb(),
		.d(n3661), .sdi(n2405), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__24__slave ( .q(_RegFile_2__24), .qb(n2406), .d(_RegFile_reg_2__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__25__master ( .q(_RegFile_reg_2__25__m2s), .qb(),
		.d(n3662), .sdi(n2406), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__25__slave ( .q(_RegFile_2__25), .qb(n2407), .d(_RegFile_reg_2__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__26__master ( .q(_RegFile_reg_2__26__m2s), .qb(),
		.d(n3663), .sdi(n2407), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__26__slave ( .q(_RegFile_2__26), .qb(n2408), .d(_RegFile_reg_2__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__27__master ( .q(_RegFile_reg_2__27__m2s), .qb(),
		.d(n3664), .sdi(n2408), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__27__slave ( .q(_RegFile_2__27), .qb(n2409), .d(_RegFile_reg_2__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__28__master ( .q(_RegFile_reg_2__28__m2s), .qb(),
		.d(n3665), .sdi(n2409), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__28__slave ( .q(_RegFile_2__28), .qb(n2410), .d(_RegFile_reg_2__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__29__master ( .q(_RegFile_reg_2__29__m2s), .qb(),
		.d(n3666), .sdi(n2410), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__29__slave ( .q(_RegFile_2__29), .qb(n2411), .d(_RegFile_reg_2__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__2__master ( .q(_RegFile_reg_2__2__m2s), .qb(),
		.d(n3639), .sdi(n4351), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n973),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__2__slave ( .q(_RegFile_2__2), .qb(n4350), .d(_RegFile_reg_2__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n973), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__30__master ( .q(_RegFile_reg_2__30__m2s), .qb(),
		.d(n3667), .sdi(n2411), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__30__slave ( .q(_RegFile_2__30), .qb(n2412), .d(_RegFile_reg_2__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__31__master ( .q(_RegFile_reg_2__31__m2s), .qb(),
		.d(n3668), .sdi(n2412), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__31__slave ( .q(_RegFile_2__31), .qb(n2413), .d(_RegFile_reg_2__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__3__master ( .q(_RegFile_reg_2__3__m2s), .qb(),
		.d(n3640), .sdi(n4350), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__3__slave ( .q(_RegFile_2__3), .qb(n4349), .d(_RegFile_reg_2__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__4__master ( .q(_RegFile_reg_2__4__m2s), .qb(),
		.d(n3641), .sdi(n4349), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__4__slave ( .q(_RegFile_2__4), .qb(n4348), .d(_RegFile_reg_2__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__5__master ( .q(_RegFile_reg_2__5__m2s), .qb(),
		.d(n3642), .sdi(n4348), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__5__slave ( .q(_RegFile_2__5), .qb(n4347), .d(_RegFile_reg_2__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__6__master ( .q(_RegFile_reg_2__6__m2s), .qb(),
		.d(n3643), .sdi(n4347), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__6__slave ( .q(_RegFile_2__6), .qb(n4346), .d(_RegFile_reg_2__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__7__master ( .q(_RegFile_reg_2__7__m2s), .qb(),
		.d(n3644), .sdi(n4346), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__7__slave ( .q(_RegFile_2__7), .qb(n4345), .d(_RegFile_reg_2__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__8__master ( .q(_RegFile_reg_2__8__m2s), .qb(),
		.d(n3645), .sdi(n4345), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__8__slave ( .q(_RegFile_2__8), .qb(n2414), .d(_RegFile_reg_2__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_2__9__master ( .q(_RegFile_reg_2__9__m2s), .qb(),
		.d(n3646), .sdi(n2414), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_2__9__slave ( .q(_RegFile_2__9), .qb(n2415), .d(_RegFile_reg_2__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__0__master ( .q(_RegFile_reg_30__0__m2s), .qb(),
		.d(n2741), .sdi(n2389), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__0__slave ( .q(_RegFile_30__0), .qb(n4128), .d(_RegFile_reg_30__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__10__master ( .q(_RegFile_reg_30__10__m2s), .qb(),
		.d(n2751), .sdi(n2439), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__10__slave ( .q(_RegFile_30__10), .qb(n2416),
		.d(_RegFile_reg_30__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__11__master ( .q(_RegFile_reg_30__11__m2s), .qb(),
		.d(n2752), .sdi(n2416), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__11__slave ( .q(_RegFile_30__11), .qb(n2417),
		.d(_RegFile_reg_30__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__12__master ( .q(_RegFile_reg_30__12__m2s), .qb(),
		.d(n2753), .sdi(n2417), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__12__slave ( .q(_RegFile_30__12), .qb(n2418),
		.d(_RegFile_reg_30__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__13__master ( .q(_RegFile_reg_30__13__m2s), .qb(),
		.d(n2754), .sdi(n2418), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__13__slave ( .q(_RegFile_30__13), .qb(n2419),
		.d(_RegFile_reg_30__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__14__master ( .q(_RegFile_reg_30__14__m2s), .qb(),
		.d(n2755), .sdi(n2419), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__14__slave ( .q(_RegFile_30__14), .qb(n2420),
		.d(_RegFile_reg_30__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__15__master ( .q(_RegFile_reg_30__15__m2s), .qb(),
		.d(n2756), .sdi(n2420), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__15__slave ( .q(_RegFile_30__15), .qb(n2421),
		.d(_RegFile_reg_30__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__16__master ( .q(_RegFile_reg_30__16__m2s), .qb(),
		.d(n2757), .sdi(n2421), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__16__slave ( .q(_RegFile_30__16), .qb(n2422),
		.d(_RegFile_reg_30__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__17__master ( .q(_RegFile_reg_30__17__m2s), .qb(),
		.d(n2758), .sdi(n2422), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__17__slave ( .q(_RegFile_30__17), .qb(n2423),
		.d(_RegFile_reg_30__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__18__master ( .q(_RegFile_reg_30__18__m2s), .qb(),
		.d(n2759), .sdi(n2423), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__18__slave ( .q(_RegFile_30__18), .qb(n2424),
		.d(_RegFile_reg_30__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__19__master ( .q(_RegFile_reg_30__19__m2s), .qb(),
		.d(n2760), .sdi(n2424), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__19__slave ( .q(_RegFile_30__19), .qb(n2425),
		.d(_RegFile_reg_30__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__1__master ( .q(_RegFile_reg_30__1__m2s), .qb(),
		.d(n2742), .sdi(n4128), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n929),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__1__slave ( .q(_RegFile_30__1), .qb(n4127), .d(_RegFile_reg_30__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n929), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__20__master ( .q(_RegFile_reg_30__20__m2s), .qb(),
		.d(n2761), .sdi(n2425), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__20__slave ( .q(_RegFile_30__20), .qb(n2426),
		.d(_RegFile_reg_30__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__21__master ( .q(_RegFile_reg_30__21__m2s), .qb(),
		.d(n2762), .sdi(n2426), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__21__slave ( .q(_RegFile_30__21), .qb(n2427),
		.d(_RegFile_reg_30__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__22__master ( .q(_RegFile_reg_30__22__m2s), .qb(),
		.d(n2763), .sdi(n2427), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__22__slave ( .q(_RegFile_30__22), .qb(n2428),
		.d(_RegFile_reg_30__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__23__master ( .q(_RegFile_reg_30__23__m2s), .qb(),
		.d(n2764), .sdi(n2428), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__23__slave ( .q(_RegFile_30__23), .qb(n2429),
		.d(_RegFile_reg_30__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__24__master ( .q(_RegFile_reg_30__24__m2s), .qb(),
		.d(n2765), .sdi(n2429), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__24__slave ( .q(_RegFile_30__24), .qb(n2430),
		.d(_RegFile_reg_30__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__25__master ( .q(_RegFile_reg_30__25__m2s), .qb(),
		.d(n2766), .sdi(n2430), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__25__slave ( .q(_RegFile_30__25), .qb(n2431),
		.d(_RegFile_reg_30__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__26__master ( .q(_RegFile_reg_30__26__m2s), .qb(),
		.d(n2767), .sdi(n2431), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__26__slave ( .q(_RegFile_30__26), .qb(n2432),
		.d(_RegFile_reg_30__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__27__master ( .q(_RegFile_reg_30__27__m2s), .qb(),
		.d(n2768), .sdi(n2432), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__27__slave ( .q(_RegFile_30__27), .qb(n2433),
		.d(_RegFile_reg_30__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__28__master ( .q(_RegFile_reg_30__28__m2s), .qb(),
		.d(n2769), .sdi(n2433), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__28__slave ( .q(_RegFile_30__28), .qb(n2434),
		.d(_RegFile_reg_30__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__29__master ( .q(_RegFile_reg_30__29__m2s), .qb(),
		.d(n2770), .sdi(n2434), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__29__slave ( .q(_RegFile_30__29), .qb(n2435),
		.d(_RegFile_reg_30__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__2__master ( .q(_RegFile_reg_30__2__m2s), .qb(),
		.d(n2743), .sdi(n4127), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n947),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__2__slave ( .q(_RegFile_30__2), .qb(n4126), .d(_RegFile_reg_30__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n947), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__30__master ( .q(_RegFile_reg_30__30__m2s), .qb(),
		.d(n2771), .sdi(n2435), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__30__slave ( .q(_RegFile_30__30), .qb(n2436),
		.d(_RegFile_reg_30__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__31__master ( .q(_RegFile_reg_30__31__m2s), .qb(),
		.d(n2772), .sdi(n2436), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__31__slave ( .q(_RegFile_30__31), .qb(n2437),
		.d(_RegFile_reg_30__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__3__master ( .q(_RegFile_reg_30__3__m2s), .qb(),
		.d(n2744), .sdi(n4126), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__3__slave ( .q(_RegFile_30__3), .qb(n4125), .d(_RegFile_reg_30__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__4__master ( .q(_RegFile_reg_30__4__m2s), .qb(),
		.d(n2745), .sdi(n4125), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__4__slave ( .q(_RegFile_30__4), .qb(n4124), .d(_RegFile_reg_30__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__5__master ( .q(_RegFile_reg_30__5__m2s), .qb(),
		.d(n2746), .sdi(n4124), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__5__slave ( .q(_RegFile_30__5), .qb(n4123), .d(_RegFile_reg_30__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__6__master ( .q(_RegFile_reg_30__6__m2s), .qb(),
		.d(n2747), .sdi(n4123), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__6__slave ( .q(_RegFile_30__6), .qb(n4122), .d(_RegFile_reg_30__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__7__master ( .q(_RegFile_reg_30__7__m2s), .qb(),
		.d(n2748), .sdi(n4122), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__7__slave ( .q(_RegFile_30__7), .qb(n4121), .d(_RegFile_reg_30__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__8__master ( .q(_RegFile_reg_30__8__m2s), .qb(),
		.d(n2749), .sdi(n4121), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__8__slave ( .q(_RegFile_30__8), .qb(n2438), .d(_RegFile_reg_30__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_30__9__master ( .q(_RegFile_reg_30__9__m2s), .qb(),
		.d(n2750), .sdi(n2438), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_30__9__slave ( .q(_RegFile_30__9), .qb(n2439), .d(_RegFile_reg_30__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__0__master ( .q(_RegFile_reg_31__0__m2s), .qb(),
		.d(n2709), .sdi(n2437), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__0__slave ( .q(_RegFile_31__0), .qb(n4120), .d(_RegFile_reg_31__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__10__master ( .q(_RegFile_reg_31__10__m2s), .qb(),
		.d(n2719), .sdi(n2463), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__10__slave ( .q(_RegFile_31__10), .qb(n2440),
		.d(_RegFile_reg_31__10__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__11__master ( .q(_RegFile_reg_31__11__m2s), .qb(),
		.d(n2720), .sdi(n2440), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__11__slave ( .q(_RegFile_31__11), .qb(n2441),
		.d(_RegFile_reg_31__11__m2s), .g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__12__master ( .q(_RegFile_reg_31__12__m2s), .qb(),
		.d(n2721), .sdi(n2441), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__12__slave ( .q(_RegFile_31__12), .qb(n2442),
		.d(_RegFile_reg_31__12__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__13__master ( .q(_RegFile_reg_31__13__m2s), .qb(),
		.d(n2722), .sdi(n2442), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__13__slave ( .q(_RegFile_31__13), .qb(n2443),
		.d(_RegFile_reg_31__13__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__14__master ( .q(_RegFile_reg_31__14__m2s), .qb(),
		.d(n2723), .sdi(n2443), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__14__slave ( .q(_RegFile_31__14), .qb(n2444),
		.d(_RegFile_reg_31__14__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__15__master ( .q(_RegFile_reg_31__15__m2s), .qb(),
		.d(n2724), .sdi(n2444), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__15__slave ( .q(_RegFile_31__15), .qb(n2445),
		.d(_RegFile_reg_31__15__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__16__master ( .q(_RegFile_reg_31__16__m2s), .qb(),
		.d(n2725), .sdi(n2445), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__16__slave ( .q(_RegFile_31__16), .qb(n2446),
		.d(_RegFile_reg_31__16__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__17__master ( .q(_RegFile_reg_31__17__m2s), .qb(),
		.d(n2726), .sdi(n2446), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__17__slave ( .q(_RegFile_31__17), .qb(n2447),
		.d(_RegFile_reg_31__17__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__18__master ( .q(_RegFile_reg_31__18__m2s), .qb(),
		.d(n2727), .sdi(n2447), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__18__slave ( .q(_RegFile_31__18), .qb(n2448),
		.d(_RegFile_reg_31__18__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__19__master ( .q(_RegFile_reg_31__19__m2s), .qb(),
		.d(n2728), .sdi(n2448), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__19__slave ( .q(_RegFile_31__19), .qb(n2449),
		.d(_RegFile_reg_31__19__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__1__master ( .q(_RegFile_reg_31__1__m2s), .qb(),
		.d(n2710), .sdi(n4120), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n928),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__1__slave ( .q(_RegFile_31__1), .qb(n4119), .d(_RegFile_reg_31__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n928), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__20__master ( .q(_RegFile_reg_31__20__m2s), .qb(),
		.d(n2729), .sdi(n2449), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__20__slave ( .q(_RegFile_31__20), .qb(n2450),
		.d(_RegFile_reg_31__20__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__21__master ( .q(_RegFile_reg_31__21__m2s), .qb(),
		.d(n2730), .sdi(n2450), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__21__slave ( .q(_RegFile_31__21), .qb(n2451),
		.d(_RegFile_reg_31__21__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__22__master ( .q(_RegFile_reg_31__22__m2s), .qb(),
		.d(n2731), .sdi(n2451), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__22__slave ( .q(_RegFile_31__22), .qb(n2452),
		.d(_RegFile_reg_31__22__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__23__master ( .q(_RegFile_reg_31__23__m2s), .qb(),
		.d(n2732), .sdi(n2452), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__23__slave ( .q(_RegFile_31__23), .qb(n2453),
		.d(_RegFile_reg_31__23__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__24__master ( .q(_RegFile_reg_31__24__m2s), .qb(),
		.d(n2733), .sdi(n2453), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__24__slave ( .q(_RegFile_31__24), .qb(n2454),
		.d(_RegFile_reg_31__24__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__25__master ( .q(_RegFile_reg_31__25__m2s), .qb(),
		.d(n2734), .sdi(n2454), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__25__slave ( .q(_RegFile_31__25), .qb(n2455),
		.d(_RegFile_reg_31__25__m2s), .g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__26__master ( .q(_RegFile_reg_31__26__m2s), .qb(),
		.d(n2735), .sdi(n2455), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__26__slave ( .q(_RegFile_31__26), .qb(n2456),
		.d(_RegFile_reg_31__26__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__27__master ( .q(_RegFile_reg_31__27__m2s), .qb(),
		.d(n2736), .sdi(n2456), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__27__slave ( .q(_RegFile_31__27), .qb(n2457),
		.d(_RegFile_reg_31__27__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__28__master ( .q(_RegFile_reg_31__28__m2s), .qb(),
		.d(n2737), .sdi(n2457), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__28__slave ( .q(_RegFile_31__28), .qb(n2458),
		.d(_RegFile_reg_31__28__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__29__master ( .q(_RegFile_reg_31__29__m2s), .qb(),
		.d(n2738), .sdi(n2458), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__29__slave ( .q(_RegFile_31__29), .qb(n2459),
		.d(_RegFile_reg_31__29__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__2__master ( .q(_RegFile_reg_31__2__m2s), .qb(),
		.d(n2711), .sdi(n4119), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n974),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__2__slave ( .q(_RegFile_31__2), .qb(n4118), .d(_RegFile_reg_31__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n974), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__30__master ( .q(_RegFile_reg_31__30__m2s), .qb(),
		.d(n2739), .sdi(n2459), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__30__slave ( .q(_RegFile_31__30), .qb(n2460),
		.d(_RegFile_reg_31__30__m2s), .g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__31__master ( .q(_RegFile_reg_31__31__m2s), .qb(),
		.d(n2740), .sdi(n2460), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__31__slave ( .q(_RegFile_31__31), .qb(n2461),
		.d(_RegFile_reg_31__31__m2s), .g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__3__master ( .q(_RegFile_reg_31__3__m2s), .qb(),
		.d(n2712), .sdi(n4118), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__3__slave ( .q(_RegFile_31__3), .qb(n4117), .d(_RegFile_reg_31__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__4__master ( .q(_RegFile_reg_31__4__m2s), .qb(),
		.d(n2713), .sdi(n4117), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__4__slave ( .q(_RegFile_31__4), .qb(n4116), .d(_RegFile_reg_31__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__5__master ( .q(_RegFile_reg_31__5__m2s), .qb(),
		.d(n2714), .sdi(n4116), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__5__slave ( .q(_RegFile_31__5), .qb(n4115), .d(_RegFile_reg_31__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__6__master ( .q(_RegFile_reg_31__6__m2s), .qb(),
		.d(n2715), .sdi(n4115), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__6__slave ( .q(_RegFile_31__6), .qb(n4114), .d(_RegFile_reg_31__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__7__master ( .q(_RegFile_reg_31__7__m2s), .qb(),
		.d(n2716), .sdi(n4114), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__7__slave ( .q(_RegFile_31__7), .qb(n4113), .d(_RegFile_reg_31__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__8__master ( .q(_RegFile_reg_31__8__m2s), .qb(),
		.d(n2717), .sdi(n4113), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__8__slave ( .q(_RegFile_31__8), .qb(n2462), .d(_RegFile_reg_31__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_31__9__master ( .q(_RegFile_reg_31__9__m2s), .qb(),
		.d(n2718), .sdi(n2462), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_31__9__slave ( .q(_RegFile_31__9), .qb(n2463), .d(_RegFile_reg_31__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__0__master ( .q(_RegFile_reg_3__0__m2s), .qb(),
		.d(n3605), .sdi(n2413), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__0__slave ( .q(_RegFile_3__0), .qb(n4344), .d(_RegFile_reg_3__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__10__master ( .q(_RegFile_reg_3__10__m2s), .qb(),
		.d(n3615), .sdi(n2487), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__10__slave ( .q(_RegFile_3__10), .qb(n2464), .d(_RegFile_reg_3__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__11__master ( .q(_RegFile_reg_3__11__m2s), .qb(),
		.d(n3616), .sdi(n2464), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__11__slave ( .q(_RegFile_3__11), .qb(n2465), .d(_RegFile_reg_3__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__12__master ( .q(_RegFile_reg_3__12__m2s), .qb(),
		.d(n3617), .sdi(n2465), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__12__slave ( .q(_RegFile_3__12), .qb(n2466), .d(_RegFile_reg_3__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__13__master ( .q(_RegFile_reg_3__13__m2s), .qb(),
		.d(n3618), .sdi(n2466), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__13__slave ( .q(_RegFile_3__13), .qb(n2467), .d(_RegFile_reg_3__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__14__master ( .q(_RegFile_reg_3__14__m2s), .qb(),
		.d(n3619), .sdi(n2467), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__14__slave ( .q(_RegFile_3__14), .qb(n2468), .d(_RegFile_reg_3__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__15__master ( .q(_RegFile_reg_3__15__m2s), .qb(),
		.d(n3620), .sdi(n2468), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__15__slave ( .q(_RegFile_3__15), .qb(n2469), .d(_RegFile_reg_3__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__16__master ( .q(_RegFile_reg_3__16__m2s), .qb(),
		.d(n3621), .sdi(n2469), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__16__slave ( .q(_RegFile_3__16), .qb(n2470), .d(_RegFile_reg_3__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__17__master ( .q(_RegFile_reg_3__17__m2s), .qb(),
		.d(n3622), .sdi(n2470), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__17__slave ( .q(_RegFile_3__17), .qb(n2471), .d(_RegFile_reg_3__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__18__master ( .q(_RegFile_reg_3__18__m2s), .qb(),
		.d(n3623), .sdi(n2471), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__18__slave ( .q(_RegFile_3__18), .qb(n2472), .d(_RegFile_reg_3__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__19__master ( .q(_RegFile_reg_3__19__m2s), .qb(),
		.d(n3624), .sdi(n2472), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__19__slave ( .q(_RegFile_3__19), .qb(n2473), .d(_RegFile_reg_3__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__1__master ( .q(_RegFile_reg_3__1__m2s), .qb(),
		.d(n3606), .sdi(n4344), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n927),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__1__slave ( .q(_RegFile_3__1), .qb(n4343), .d(_RegFile_reg_3__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n927), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__20__master ( .q(_RegFile_reg_3__20__m2s), .qb(),
		.d(n3625), .sdi(n2473), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__20__slave ( .q(_RegFile_3__20), .qb(n2474), .d(_RegFile_reg_3__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__21__master ( .q(_RegFile_reg_3__21__m2s), .qb(),
		.d(n3626), .sdi(n2474), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__21__slave ( .q(_RegFile_3__21), .qb(n2475), .d(_RegFile_reg_3__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__22__master ( .q(_RegFile_reg_3__22__m2s), .qb(),
		.d(n3627), .sdi(n2475), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__22__slave ( .q(_RegFile_3__22), .qb(n2476), .d(_RegFile_reg_3__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__23__master ( .q(_RegFile_reg_3__23__m2s), .qb(),
		.d(n3628), .sdi(n2476), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__23__slave ( .q(_RegFile_3__23), .qb(n2477), .d(_RegFile_reg_3__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__24__master ( .q(_RegFile_reg_3__24__m2s), .qb(),
		.d(n3629), .sdi(n2477), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__24__slave ( .q(_RegFile_3__24), .qb(n2478), .d(_RegFile_reg_3__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__25__master ( .q(_RegFile_reg_3__25__m2s), .qb(),
		.d(n3630), .sdi(n2478), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__25__slave ( .q(_RegFile_3__25), .qb(n2479), .d(_RegFile_reg_3__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__26__master ( .q(_RegFile_reg_3__26__m2s), .qb(),
		.d(n3631), .sdi(n2479), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__26__slave ( .q(_RegFile_3__26), .qb(n2480), .d(_RegFile_reg_3__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__27__master ( .q(_RegFile_reg_3__27__m2s), .qb(),
		.d(n3632), .sdi(n2480), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__27__slave ( .q(_RegFile_3__27), .qb(n2481), .d(_RegFile_reg_3__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__28__master ( .q(_RegFile_reg_3__28__m2s), .qb(),
		.d(n3633), .sdi(n2481), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__28__slave ( .q(_RegFile_3__28), .qb(n2482), .d(_RegFile_reg_3__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__29__master ( .q(_RegFile_reg_3__29__m2s), .qb(),
		.d(n3634), .sdi(n2482), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__29__slave ( .q(_RegFile_3__29), .qb(n2483), .d(_RegFile_reg_3__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__2__master ( .q(_RegFile_reg_3__2__m2s), .qb(),
		.d(n3607), .sdi(n4343), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n975),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__2__slave ( .q(_RegFile_3__2), .qb(n4342), .d(_RegFile_reg_3__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n975), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__30__master ( .q(_RegFile_reg_3__30__m2s), .qb(),
		.d(n3635), .sdi(n2483), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__30__slave ( .q(_RegFile_3__30), .qb(n2484), .d(_RegFile_reg_3__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__31__master ( .q(_RegFile_reg_3__31__m2s), .qb(),
		.d(n3636), .sdi(n2484), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__31__slave ( .q(_RegFile_3__31), .qb(n2485), .d(_RegFile_reg_3__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__3__master ( .q(_RegFile_reg_3__3__m2s), .qb(),
		.d(n3608), .sdi(n4342), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__3__slave ( .q(_RegFile_3__3), .qb(n4341), .d(_RegFile_reg_3__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__4__master ( .q(_RegFile_reg_3__4__m2s), .qb(),
		.d(n3609), .sdi(n4341), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__4__slave ( .q(_RegFile_3__4), .qb(n4340), .d(_RegFile_reg_3__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__5__master ( .q(_RegFile_reg_3__5__m2s), .qb(),
		.d(n3610), .sdi(n4340), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__5__slave ( .q(_RegFile_3__5), .qb(n4339), .d(_RegFile_reg_3__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__6__master ( .q(_RegFile_reg_3__6__m2s), .qb(),
		.d(n3611), .sdi(n4339), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__6__slave ( .q(_RegFile_3__6), .qb(n4338), .d(_RegFile_reg_3__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__7__master ( .q(_RegFile_reg_3__7__m2s), .qb(),
		.d(n3612), .sdi(n4338), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__7__slave ( .q(_RegFile_3__7), .qb(n4337), .d(_RegFile_reg_3__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__8__master ( .q(_RegFile_reg_3__8__m2s), .qb(),
		.d(n3613), .sdi(n4337), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__8__slave ( .q(_RegFile_3__8), .qb(n2486), .d(_RegFile_reg_3__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_3__9__master ( .q(_RegFile_reg_3__9__m2s), .qb(),
		.d(n3614), .sdi(n2486), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n926),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_3__9__slave ( .q(_RegFile_3__9), .qb(n2487), .d(_RegFile_reg_3__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n926), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__0__master ( .q(_RegFile_reg_4__0__m2s), .qb(),
		.d(n3573), .sdi(n2485), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__0__slave ( .q(_RegFile_4__0), .qb(n4336), .d(_RegFile_reg_4__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__10__master ( .q(_RegFile_reg_4__10__m2s), .qb(),
		.d(n3583), .sdi(n2511), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__10__slave ( .q(_RegFile_4__10), .qb(n2488), .d(_RegFile_reg_4__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__11__master ( .q(_RegFile_reg_4__11__m2s), .qb(),
		.d(n3584), .sdi(n2488), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__11__slave ( .q(_RegFile_4__11), .qb(n2489), .d(_RegFile_reg_4__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__12__master ( .q(_RegFile_reg_4__12__m2s), .qb(),
		.d(n3585), .sdi(n2489), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__12__slave ( .q(_RegFile_4__12), .qb(n2490), .d(_RegFile_reg_4__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__13__master ( .q(_RegFile_reg_4__13__m2s), .qb(),
		.d(n3586), .sdi(n2490), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__13__slave ( .q(_RegFile_4__13), .qb(n2491), .d(_RegFile_reg_4__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__14__master ( .q(_RegFile_reg_4__14__m2s), .qb(),
		.d(n3587), .sdi(n2491), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__14__slave ( .q(_RegFile_4__14), .qb(n2492), .d(_RegFile_reg_4__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__15__master ( .q(_RegFile_reg_4__15__m2s), .qb(),
		.d(n3588), .sdi(n2492), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__15__slave ( .q(_RegFile_4__15), .qb(n2493), .d(_RegFile_reg_4__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__16__master ( .q(_RegFile_reg_4__16__m2s), .qb(),
		.d(n3589), .sdi(n2493), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__16__slave ( .q(_RegFile_4__16), .qb(n2494), .d(_RegFile_reg_4__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__17__master ( .q(_RegFile_reg_4__17__m2s), .qb(),
		.d(n3590), .sdi(n2494), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__17__slave ( .q(_RegFile_4__17), .qb(n2495), .d(_RegFile_reg_4__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__18__master ( .q(_RegFile_reg_4__18__m2s), .qb(),
		.d(n3591), .sdi(n2495), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__18__slave ( .q(_RegFile_4__18), .qb(n2496), .d(_RegFile_reg_4__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__19__master ( .q(_RegFile_reg_4__19__m2s), .qb(),
		.d(n3592), .sdi(n2496), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__19__slave ( .q(_RegFile_4__19), .qb(n2497), .d(_RegFile_reg_4__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__1__master ( .q(_RegFile_reg_4__1__m2s), .qb(),
		.d(n3574), .sdi(n4336), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__1__slave ( .q(_RegFile_4__1), .qb(n4335), .d(_RegFile_reg_4__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__20__master ( .q(_RegFile_reg_4__20__m2s), .qb(),
		.d(n3593), .sdi(n2497), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__20__slave ( .q(_RegFile_4__20), .qb(n2498), .d(_RegFile_reg_4__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__21__master ( .q(_RegFile_reg_4__21__m2s), .qb(),
		.d(n3594), .sdi(n2498), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__21__slave ( .q(_RegFile_4__21), .qb(n2499), .d(_RegFile_reg_4__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__22__master ( .q(_RegFile_reg_4__22__m2s), .qb(),
		.d(n3595), .sdi(n2499), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__22__slave ( .q(_RegFile_4__22), .qb(n2500), .d(_RegFile_reg_4__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__23__master ( .q(_RegFile_reg_4__23__m2s), .qb(),
		.d(n3596), .sdi(n2500), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__23__slave ( .q(_RegFile_4__23), .qb(n2501), .d(_RegFile_reg_4__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__24__master ( .q(_RegFile_reg_4__24__m2s), .qb(),
		.d(n3597), .sdi(n2501), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__24__slave ( .q(_RegFile_4__24), .qb(n2502), .d(_RegFile_reg_4__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__25__master ( .q(_RegFile_reg_4__25__m2s), .qb(),
		.d(n3598), .sdi(n2502), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__25__slave ( .q(_RegFile_4__25), .qb(n2503), .d(_RegFile_reg_4__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__26__master ( .q(_RegFile_reg_4__26__m2s), .qb(),
		.d(n3599), .sdi(n2503), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__26__slave ( .q(_RegFile_4__26), .qb(n2504), .d(_RegFile_reg_4__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__27__master ( .q(_RegFile_reg_4__27__m2s), .qb(),
		.d(n3600), .sdi(n2504), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__27__slave ( .q(_RegFile_4__27), .qb(n2505), .d(_RegFile_reg_4__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__28__master ( .q(_RegFile_reg_4__28__m2s), .qb(),
		.d(n3601), .sdi(n2505), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__28__slave ( .q(_RegFile_4__28), .qb(n2506), .d(_RegFile_reg_4__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__29__master ( .q(_RegFile_reg_4__29__m2s), .qb(),
		.d(n3602), .sdi(n2506), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__29__slave ( .q(_RegFile_4__29), .qb(n2507), .d(_RegFile_reg_4__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__2__master ( .q(_RegFile_reg_4__2__m2s), .qb(),
		.d(n3575), .sdi(n4335), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n976),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__2__slave ( .q(_RegFile_4__2), .qb(n4334), .d(_RegFile_reg_4__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n976), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__30__master ( .q(_RegFile_reg_4__30__m2s), .qb(),
		.d(n3603), .sdi(n2507), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__30__slave ( .q(_RegFile_4__30), .qb(n2508), .d(_RegFile_reg_4__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__31__master ( .q(_RegFile_reg_4__31__m2s), .qb(),
		.d(n3604), .sdi(n2508), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__31__slave ( .q(_RegFile_4__31), .qb(n2509), .d(_RegFile_reg_4__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__3__master ( .q(_RegFile_reg_4__3__m2s), .qb(),
		.d(n3576), .sdi(n4334), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__3__slave ( .q(_RegFile_4__3), .qb(n4333), .d(_RegFile_reg_4__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__4__master ( .q(_RegFile_reg_4__4__m2s), .qb(),
		.d(n3577), .sdi(n4333), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__4__slave ( .q(_RegFile_4__4), .qb(n4332), .d(_RegFile_reg_4__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__5__master ( .q(_RegFile_reg_4__5__m2s), .qb(),
		.d(n3578), .sdi(n4332), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__5__slave ( .q(_RegFile_4__5), .qb(n4331), .d(_RegFile_reg_4__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__6__master ( .q(_RegFile_reg_4__6__m2s), .qb(),
		.d(n3579), .sdi(n4331), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__6__slave ( .q(_RegFile_4__6), .qb(n4330), .d(_RegFile_reg_4__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__7__master ( .q(_RegFile_reg_4__7__m2s), .qb(),
		.d(n3580), .sdi(n4330), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n925),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__7__slave ( .q(_RegFile_4__7), .qb(n4329), .d(_RegFile_reg_4__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n925), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__8__master ( .q(_RegFile_reg_4__8__m2s), .qb(),
		.d(n3581), .sdi(n4329), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__8__slave ( .q(_RegFile_4__8), .qb(n2510), .d(_RegFile_reg_4__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_4__9__master ( .q(_RegFile_reg_4__9__m2s), .qb(),
		.d(n3582), .sdi(n2510), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_4__9__slave ( .q(_RegFile_4__9), .qb(n2511), .d(_RegFile_reg_4__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__0__master ( .q(_RegFile_reg_5__0__m2s), .qb(),
		.d(n3541), .sdi(n2509), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__0__slave ( .q(_RegFile_5__0), .qb(n4328), .d(_RegFile_reg_5__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__10__master ( .q(_RegFile_reg_5__10__m2s), .qb(),
		.d(n3551), .sdi(n2535), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__10__slave ( .q(_RegFile_5__10), .qb(n2512), .d(_RegFile_reg_5__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__11__master ( .q(_RegFile_reg_5__11__m2s), .qb(),
		.d(n3552), .sdi(n2512), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__11__slave ( .q(_RegFile_5__11), .qb(n2513), .d(_RegFile_reg_5__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__12__master ( .q(_RegFile_reg_5__12__m2s), .qb(),
		.d(n3553), .sdi(n2513), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__12__slave ( .q(_RegFile_5__12), .qb(n2514), .d(_RegFile_reg_5__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__13__master ( .q(_RegFile_reg_5__13__m2s), .qb(),
		.d(n3554), .sdi(n2514), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__13__slave ( .q(_RegFile_5__13), .qb(n2515), .d(_RegFile_reg_5__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__14__master ( .q(_RegFile_reg_5__14__m2s), .qb(),
		.d(n3555), .sdi(n2515), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__14__slave ( .q(_RegFile_5__14), .qb(n2516), .d(_RegFile_reg_5__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__15__master ( .q(_RegFile_reg_5__15__m2s), .qb(),
		.d(n3556), .sdi(n2516), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__15__slave ( .q(_RegFile_5__15), .qb(n2517), .d(_RegFile_reg_5__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__16__master ( .q(_RegFile_reg_5__16__m2s), .qb(),
		.d(n3557), .sdi(n2517), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__16__slave ( .q(_RegFile_5__16), .qb(n2518), .d(_RegFile_reg_5__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__17__master ( .q(_RegFile_reg_5__17__m2s), .qb(),
		.d(n3558), .sdi(n2518), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__17__slave ( .q(_RegFile_5__17), .qb(n2519), .d(_RegFile_reg_5__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__18__master ( .q(_RegFile_reg_5__18__m2s), .qb(),
		.d(n3559), .sdi(n2519), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__18__slave ( .q(_RegFile_5__18), .qb(n2520), .d(_RegFile_reg_5__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__19__master ( .q(_RegFile_reg_5__19__m2s), .qb(),
		.d(n3560), .sdi(n2520), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__19__slave ( .q(_RegFile_5__19), .qb(n2521), .d(_RegFile_reg_5__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__1__master ( .q(_RegFile_reg_5__1__m2s), .qb(),
		.d(n3542), .sdi(n4328), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__1__slave ( .q(_RegFile_5__1), .qb(n4327), .d(_RegFile_reg_5__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__20__master ( .q(_RegFile_reg_5__20__m2s), .qb(),
		.d(n3561), .sdi(n2521), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__20__slave ( .q(_RegFile_5__20), .qb(n2522), .d(_RegFile_reg_5__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__21__master ( .q(_RegFile_reg_5__21__m2s), .qb(),
		.d(n3562), .sdi(n2522), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__21__slave ( .q(_RegFile_5__21), .qb(n2523), .d(_RegFile_reg_5__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__22__master ( .q(_RegFile_reg_5__22__m2s), .qb(),
		.d(n3563), .sdi(n2523), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__22__slave ( .q(_RegFile_5__22), .qb(n2524), .d(_RegFile_reg_5__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__23__master ( .q(_RegFile_reg_5__23__m2s), .qb(),
		.d(n3564), .sdi(n2524), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__23__slave ( .q(_RegFile_5__23), .qb(n2525), .d(_RegFile_reg_5__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__24__master ( .q(_RegFile_reg_5__24__m2s), .qb(),
		.d(n3565), .sdi(n2525), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__24__slave ( .q(_RegFile_5__24), .qb(n2526), .d(_RegFile_reg_5__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__25__master ( .q(_RegFile_reg_5__25__m2s), .qb(),
		.d(n3566), .sdi(n2526), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__25__slave ( .q(_RegFile_5__25), .qb(n2527), .d(_RegFile_reg_5__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__26__master ( .q(_RegFile_reg_5__26__m2s), .qb(),
		.d(n3567), .sdi(n2527), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__26__slave ( .q(_RegFile_5__26), .qb(n2528), .d(_RegFile_reg_5__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__27__master ( .q(_RegFile_reg_5__27__m2s), .qb(),
		.d(n3568), .sdi(n2528), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__27__slave ( .q(_RegFile_5__27), .qb(n2529), .d(_RegFile_reg_5__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__28__master ( .q(_RegFile_reg_5__28__m2s), .qb(),
		.d(n3569), .sdi(n2529), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__28__slave ( .q(_RegFile_5__28), .qb(n2530), .d(_RegFile_reg_5__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__29__master ( .q(_RegFile_reg_5__29__m2s), .qb(),
		.d(n3570), .sdi(n2530), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__29__slave ( .q(_RegFile_5__29), .qb(n2531), .d(_RegFile_reg_5__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__2__master ( .q(_RegFile_reg_5__2__m2s), .qb(),
		.d(n3543), .sdi(n4327), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n977),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__2__slave ( .q(_RegFile_5__2), .qb(n4326), .d(_RegFile_reg_5__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n977), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__30__master ( .q(_RegFile_reg_5__30__m2s), .qb(),
		.d(n3571), .sdi(n2531), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__30__slave ( .q(_RegFile_5__30), .qb(n2532), .d(_RegFile_reg_5__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__31__master ( .q(_RegFile_reg_5__31__m2s), .qb(),
		.d(n3572), .sdi(n2532), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__31__slave ( .q(_RegFile_5__31), .qb(n2533), .d(_RegFile_reg_5__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__3__master ( .q(_RegFile_reg_5__3__m2s), .qb(),
		.d(n3544), .sdi(n4326), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__3__slave ( .q(_RegFile_5__3), .qb(n4325), .d(_RegFile_reg_5__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__4__master ( .q(_RegFile_reg_5__4__m2s), .qb(),
		.d(n3545), .sdi(n4325), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__4__slave ( .q(_RegFile_5__4), .qb(n4324), .d(_RegFile_reg_5__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__5__master ( .q(_RegFile_reg_5__5__m2s), .qb(),
		.d(n3546), .sdi(n4324), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n924),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__5__slave ( .q(_RegFile_5__5), .qb(n4323), .d(_RegFile_reg_5__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n924), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__6__master ( .q(_RegFile_reg_5__6__m2s), .qb(),
		.d(n3547), .sdi(n4323), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__6__slave ( .q(_RegFile_5__6), .qb(n4322), .d(_RegFile_reg_5__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__7__master ( .q(_RegFile_reg_5__7__m2s), .qb(),
		.d(n3548), .sdi(n4322), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__7__slave ( .q(_RegFile_5__7), .qb(n4321), .d(_RegFile_reg_5__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__8__master ( .q(_RegFile_reg_5__8__m2s), .qb(),
		.d(n3549), .sdi(n4321), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__8__slave ( .q(_RegFile_5__8), .qb(n2534), .d(_RegFile_reg_5__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_5__9__master ( .q(_RegFile_reg_5__9__m2s), .qb(),
		.d(n3550), .sdi(n2534), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_5__9__slave ( .q(_RegFile_5__9), .qb(n2535), .d(_RegFile_reg_5__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__0__master ( .q(_RegFile_reg_6__0__m2s), .qb(),
		.d(n3509), .sdi(n2533), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__0__slave ( .q(_RegFile_6__0), .qb(n4320), .d(_RegFile_reg_6__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__10__master ( .q(_RegFile_reg_6__10__m2s), .qb(),
		.d(n3519), .sdi(n2559), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__10__slave ( .q(_RegFile_6__10), .qb(n2536), .d(_RegFile_reg_6__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__11__master ( .q(_RegFile_reg_6__11__m2s), .qb(),
		.d(n3520), .sdi(n2536), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__11__slave ( .q(_RegFile_6__11), .qb(n2537), .d(_RegFile_reg_6__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__12__master ( .q(_RegFile_reg_6__12__m2s), .qb(),
		.d(n3521), .sdi(n2537), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__12__slave ( .q(_RegFile_6__12), .qb(n2538), .d(_RegFile_reg_6__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__13__master ( .q(_RegFile_reg_6__13__m2s), .qb(),
		.d(n3522), .sdi(n2538), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__13__slave ( .q(_RegFile_6__13), .qb(n2539), .d(_RegFile_reg_6__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__14__master ( .q(_RegFile_reg_6__14__m2s), .qb(),
		.d(n3523), .sdi(n2539), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__14__slave ( .q(_RegFile_6__14), .qb(n2540), .d(_RegFile_reg_6__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__15__master ( .q(_RegFile_reg_6__15__m2s), .qb(),
		.d(n3524), .sdi(n2540), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__15__slave ( .q(_RegFile_6__15), .qb(n2541), .d(_RegFile_reg_6__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__16__master ( .q(_RegFile_reg_6__16__m2s), .qb(),
		.d(n3525), .sdi(n2541), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__16__slave ( .q(_RegFile_6__16), .qb(n2542), .d(_RegFile_reg_6__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__17__master ( .q(_RegFile_reg_6__17__m2s), .qb(),
		.d(n3526), .sdi(n2542), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__17__slave ( .q(_RegFile_6__17), .qb(n2543), .d(_RegFile_reg_6__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__18__master ( .q(_RegFile_reg_6__18__m2s), .qb(),
		.d(n3527), .sdi(n2543), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n978),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__18__slave ( .q(_RegFile_6__18), .qb(n2544), .d(_RegFile_reg_6__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n978), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__19__master ( .q(_RegFile_reg_6__19__m2s), .qb(),
		.d(n3528), .sdi(n2544), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__19__slave ( .q(_RegFile_6__19), .qb(n2545), .d(_RegFile_reg_6__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__1__master ( .q(_RegFile_reg_6__1__m2s), .qb(),
		.d(n3510), .sdi(n4320), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__1__slave ( .q(_RegFile_6__1), .qb(n4319), .d(_RegFile_reg_6__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__20__master ( .q(_RegFile_reg_6__20__m2s), .qb(),
		.d(n3529), .sdi(n2545), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__20__slave ( .q(_RegFile_6__20), .qb(n2546), .d(_RegFile_reg_6__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__21__master ( .q(_RegFile_reg_6__21__m2s), .qb(),
		.d(n3530), .sdi(n2546), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__21__slave ( .q(_RegFile_6__21), .qb(n2547), .d(_RegFile_reg_6__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__22__master ( .q(_RegFile_reg_6__22__m2s), .qb(),
		.d(n3531), .sdi(n2547), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__22__slave ( .q(_RegFile_6__22), .qb(n2548), .d(_RegFile_reg_6__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__23__master ( .q(_RegFile_reg_6__23__m2s), .qb(),
		.d(n3532), .sdi(n2548), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__23__slave ( .q(_RegFile_6__23), .qb(n2549), .d(_RegFile_reg_6__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__24__master ( .q(_RegFile_reg_6__24__m2s), .qb(),
		.d(n3533), .sdi(n2549), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__24__slave ( .q(_RegFile_6__24), .qb(n2550), .d(_RegFile_reg_6__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__25__master ( .q(_RegFile_reg_6__25__m2s), .qb(),
		.d(n3534), .sdi(n2550), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__25__slave ( .q(_RegFile_6__25), .qb(n2551), .d(_RegFile_reg_6__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__26__master ( .q(_RegFile_reg_6__26__m2s), .qb(),
		.d(n3535), .sdi(n2551), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__26__slave ( .q(_RegFile_6__26), .qb(n2552), .d(_RegFile_reg_6__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__27__master ( .q(_RegFile_reg_6__27__m2s), .qb(),
		.d(n3536), .sdi(n2552), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__27__slave ( .q(_RegFile_6__27), .qb(n2553), .d(_RegFile_reg_6__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__28__master ( .q(_RegFile_reg_6__28__m2s), .qb(),
		.d(n3537), .sdi(n2553), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__28__slave ( .q(_RegFile_6__28), .qb(n2554), .d(_RegFile_reg_6__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__29__master ( .q(_RegFile_reg_6__29__m2s), .qb(),
		.d(n3538), .sdi(n2554), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__29__slave ( .q(_RegFile_6__29), .qb(n2555), .d(_RegFile_reg_6__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__2__master ( .q(_RegFile_reg_6__2__m2s), .qb(),
		.d(n3511), .sdi(n4319), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__2__slave ( .q(_RegFile_6__2), .qb(n4318), .d(_RegFile_reg_6__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__30__master ( .q(_RegFile_reg_6__30__m2s), .qb(),
		.d(n3539), .sdi(n2555), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__30__slave ( .q(_RegFile_6__30), .qb(n2556), .d(_RegFile_reg_6__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__31__master ( .q(_RegFile_reg_6__31__m2s), .qb(),
		.d(n3540), .sdi(n2556), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__31__slave ( .q(_RegFile_6__31), .qb(n2557), .d(_RegFile_reg_6__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__3__master ( .q(_RegFile_reg_6__3__m2s), .qb(),
		.d(n3512), .sdi(n4318), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n923),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__3__slave ( .q(_RegFile_6__3), .qb(n4317), .d(_RegFile_reg_6__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n923), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__4__master ( .q(_RegFile_reg_6__4__m2s), .qb(),
		.d(n3513), .sdi(n4317), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__4__slave ( .q(_RegFile_6__4), .qb(n4316), .d(_RegFile_reg_6__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__5__master ( .q(_RegFile_reg_6__5__m2s), .qb(),
		.d(n3514), .sdi(n4316), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__5__slave ( .q(_RegFile_6__5), .qb(n4315), .d(_RegFile_reg_6__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__6__master ( .q(_RegFile_reg_6__6__m2s), .qb(),
		.d(n3515), .sdi(n4315), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__6__slave ( .q(_RegFile_6__6), .qb(n4314), .d(_RegFile_reg_6__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__7__master ( .q(_RegFile_reg_6__7__m2s), .qb(),
		.d(n3516), .sdi(n4314), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__7__slave ( .q(_RegFile_6__7), .qb(n4313), .d(_RegFile_reg_6__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__8__master ( .q(_RegFile_reg_6__8__m2s), .qb(),
		.d(n3517), .sdi(n4313), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__8__slave ( .q(_RegFile_6__8), .qb(n2558), .d(_RegFile_reg_6__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_6__9__master ( .q(_RegFile_reg_6__9__m2s), .qb(),
		.d(n3518), .sdi(n2558), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_6__9__slave ( .q(_RegFile_6__9), .qb(n2559), .d(_RegFile_reg_6__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__0__master ( .q(_RegFile_reg_7__0__m2s), .qb(),
		.d(n3477), .sdi(n2557), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__0__slave ( .q(_RegFile_7__0), .qb(n4312), .d(_RegFile_reg_7__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__10__master ( .q(_RegFile_reg_7__10__m2s), .qb(),
		.d(n3487), .sdi(n2583), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__10__slave ( .q(_RegFile_7__10), .qb(n2560), .d(_RegFile_reg_7__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__11__master ( .q(_RegFile_reg_7__11__m2s), .qb(),
		.d(n3488), .sdi(n2560), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__11__slave ( .q(_RegFile_7__11), .qb(n2561), .d(_RegFile_reg_7__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__12__master ( .q(_RegFile_reg_7__12__m2s), .qb(),
		.d(n3489), .sdi(n2561), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__12__slave ( .q(_RegFile_7__12), .qb(n2562), .d(_RegFile_reg_7__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__13__master ( .q(_RegFile_reg_7__13__m2s), .qb(),
		.d(n3490), .sdi(n2562), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__13__slave ( .q(_RegFile_7__13), .qb(n2563), .d(_RegFile_reg_7__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__14__master ( .q(_RegFile_reg_7__14__m2s), .qb(),
		.d(n3491), .sdi(n2563), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__14__slave ( .q(_RegFile_7__14), .qb(n2564), .d(_RegFile_reg_7__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__15__master ( .q(_RegFile_reg_7__15__m2s), .qb(),
		.d(n3492), .sdi(n2564), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__15__slave ( .q(_RegFile_7__15), .qb(n2565), .d(_RegFile_reg_7__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__16__master ( .q(_RegFile_reg_7__16__m2s), .qb(),
		.d(n3493), .sdi(n2565), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n979),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__16__slave ( .q(_RegFile_7__16), .qb(n2566), .d(_RegFile_reg_7__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n979), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__17__master ( .q(_RegFile_reg_7__17__m2s), .qb(),
		.d(n3494), .sdi(n2566), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__17__slave ( .q(_RegFile_7__17), .qb(n2567), .d(_RegFile_reg_7__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__18__master ( .q(_RegFile_reg_7__18__m2s), .qb(),
		.d(n3495), .sdi(n2567), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__18__slave ( .q(_RegFile_7__18), .qb(n2568), .d(_RegFile_reg_7__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__19__master ( .q(_RegFile_reg_7__19__m2s), .qb(),
		.d(n3496), .sdi(n2568), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__19__slave ( .q(_RegFile_7__19), .qb(n2569), .d(_RegFile_reg_7__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__1__master ( .q(_RegFile_reg_7__1__m2s), .qb(),
		.d(n3478), .sdi(n4312), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__1__slave ( .q(_RegFile_7__1), .qb(n4311), .d(_RegFile_reg_7__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__20__master ( .q(_RegFile_reg_7__20__m2s), .qb(),
		.d(n3497), .sdi(n2569), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__20__slave ( .q(_RegFile_7__20), .qb(n2570), .d(_RegFile_reg_7__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__21__master ( .q(_RegFile_reg_7__21__m2s), .qb(),
		.d(n3498), .sdi(n2570), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__21__slave ( .q(_RegFile_7__21), .qb(n2571), .d(_RegFile_reg_7__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__22__master ( .q(_RegFile_reg_7__22__m2s), .qb(),
		.d(n3499), .sdi(n2571), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__22__slave ( .q(_RegFile_7__22), .qb(n2572), .d(_RegFile_reg_7__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__23__master ( .q(_RegFile_reg_7__23__m2s), .qb(),
		.d(n3500), .sdi(n2572), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__23__slave ( .q(_RegFile_7__23), .qb(n2573), .d(_RegFile_reg_7__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__24__master ( .q(_RegFile_reg_7__24__m2s), .qb(),
		.d(n3501), .sdi(n2573), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__24__slave ( .q(_RegFile_7__24), .qb(n2574), .d(_RegFile_reg_7__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__25__master ( .q(_RegFile_reg_7__25__m2s), .qb(),
		.d(n3502), .sdi(n2574), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__25__slave ( .q(_RegFile_7__25), .qb(n2575), .d(_RegFile_reg_7__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__26__master ( .q(_RegFile_reg_7__26__m2s), .qb(),
		.d(n3503), .sdi(n2575), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__26__slave ( .q(_RegFile_7__26), .qb(n2576), .d(_RegFile_reg_7__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__27__master ( .q(_RegFile_reg_7__27__m2s), .qb(),
		.d(n3504), .sdi(n2576), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__27__slave ( .q(_RegFile_7__27), .qb(n2577), .d(_RegFile_reg_7__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__28__master ( .q(_RegFile_reg_7__28__m2s), .qb(),
		.d(n3505), .sdi(n2577), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__28__slave ( .q(_RegFile_7__28), .qb(n2578), .d(_RegFile_reg_7__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__29__master ( .q(_RegFile_reg_7__29__m2s), .qb(),
		.d(n3506), .sdi(n2578), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__29__slave ( .q(_RegFile_7__29), .qb(n2579), .d(_RegFile_reg_7__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__2__master ( .q(_RegFile_reg_7__2__m2s), .qb(),
		.d(n3479), .sdi(n4311), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__2__slave ( .q(_RegFile_7__2), .qb(n4310), .d(_RegFile_reg_7__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__30__master ( .q(_RegFile_reg_7__30__m2s), .qb(),
		.d(n3507), .sdi(n2579), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__30__slave ( .q(_RegFile_7__30), .qb(n2580), .d(_RegFile_reg_7__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__31__master ( .q(_RegFile_reg_7__31__m2s), .qb(),
		.d(n3508), .sdi(n2580), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__31__slave ( .q(_RegFile_7__31), .qb(n2581), .d(_RegFile_reg_7__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__3__master ( .q(_RegFile_reg_7__3__m2s), .qb(),
		.d(n3480), .sdi(n4310), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n922),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__3__slave ( .q(_RegFile_7__3), .qb(n4309), .d(_RegFile_reg_7__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n922), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__4__master ( .q(_RegFile_reg_7__4__m2s), .qb(),
		.d(n3481), .sdi(n4309), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__4__slave ( .q(_RegFile_7__4), .qb(n4308), .d(_RegFile_reg_7__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__5__master ( .q(_RegFile_reg_7__5__m2s), .qb(),
		.d(n3482), .sdi(n4308), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__5__slave ( .q(_RegFile_7__5), .qb(n4307), .d(_RegFile_reg_7__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__6__master ( .q(_RegFile_reg_7__6__m2s), .qb(),
		.d(n3483), .sdi(n4307), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__6__slave ( .q(_RegFile_7__6), .qb(n4306), .d(_RegFile_reg_7__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__7__master ( .q(_RegFile_reg_7__7__m2s), .qb(),
		.d(n3484), .sdi(n4306), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__7__slave ( .q(_RegFile_7__7), .qb(n4305), .d(_RegFile_reg_7__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__8__master ( .q(_RegFile_reg_7__8__m2s), .qb(),
		.d(n3485), .sdi(n4305), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__8__slave ( .q(_RegFile_7__8), .qb(n2582), .d(_RegFile_reg_7__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_7__9__master ( .q(_RegFile_reg_7__9__m2s), .qb(),
		.d(n3486), .sdi(n2582), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_7__9__slave ( .q(_RegFile_7__9), .qb(n2583), .d(_RegFile_reg_7__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__0__master ( .q(_RegFile_reg_8__0__m2s), .qb(),
		.d(n3445), .sdi(n2581), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__0__slave ( .q(_RegFile_8__0), .qb(n4304), .d(_RegFile_reg_8__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__10__master ( .q(_RegFile_reg_8__10__m2s), .qb(),
		.d(n3455), .sdi(n2607), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__10__slave ( .q(_RegFile_8__10), .qb(n2584), .d(_RegFile_reg_8__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__11__master ( .q(_RegFile_reg_8__11__m2s), .qb(),
		.d(n3456), .sdi(n2584), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__11__slave ( .q(_RegFile_8__11), .qb(n2585), .d(_RegFile_reg_8__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__12__master ( .q(_RegFile_reg_8__12__m2s), .qb(),
		.d(n3457), .sdi(n2585), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__12__slave ( .q(_RegFile_8__12), .qb(n2586), .d(_RegFile_reg_8__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__13__master ( .q(_RegFile_reg_8__13__m2s), .qb(),
		.d(n3458), .sdi(n2586), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__13__slave ( .q(_RegFile_8__13), .qb(n2587), .d(_RegFile_reg_8__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__14__master ( .q(_RegFile_reg_8__14__m2s), .qb(),
		.d(n3459), .sdi(n2587), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__14__slave ( .q(_RegFile_8__14), .qb(n2588), .d(_RegFile_reg_8__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__15__master ( .q(_RegFile_reg_8__15__m2s), .qb(),
		.d(n3460), .sdi(n2588), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__15__slave ( .q(_RegFile_8__15), .qb(n2589), .d(_RegFile_reg_8__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__16__master ( .q(_RegFile_reg_8__16__m2s), .qb(),
		.d(n3461), .sdi(n2589), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__16__slave ( .q(_RegFile_8__16), .qb(n2590), .d(_RegFile_reg_8__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__17__master ( .q(_RegFile_reg_8__17__m2s), .qb(),
		.d(n3462), .sdi(n2590), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__17__slave ( .q(_RegFile_8__17), .qb(n2591), .d(_RegFile_reg_8__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__18__master ( .q(_RegFile_reg_8__18__m2s), .qb(),
		.d(n3463), .sdi(n2591), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__18__slave ( .q(_RegFile_8__18), .qb(n2592), .d(_RegFile_reg_8__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__19__master ( .q(_RegFile_reg_8__19__m2s), .qb(),
		.d(n3464), .sdi(n2592), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__19__slave ( .q(_RegFile_8__19), .qb(n2593), .d(_RegFile_reg_8__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__1__master ( .q(_RegFile_reg_8__1__m2s), .qb(),
		.d(n3446), .sdi(n4304), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__1__slave ( .q(_RegFile_8__1), .qb(n4303), .d(_RegFile_reg_8__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__20__master ( .q(_RegFile_reg_8__20__m2s), .qb(),
		.d(n3465), .sdi(n2593), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__20__slave ( .q(_RegFile_8__20), .qb(n2594), .d(_RegFile_reg_8__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__21__master ( .q(_RegFile_reg_8__21__m2s), .qb(),
		.d(n3466), .sdi(n2594), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__21__slave ( .q(_RegFile_8__21), .qb(n2595), .d(_RegFile_reg_8__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__22__master ( .q(_RegFile_reg_8__22__m2s), .qb(),
		.d(n3467), .sdi(n2595), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__22__slave ( .q(_RegFile_8__22), .qb(n2596), .d(_RegFile_reg_8__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__23__master ( .q(_RegFile_reg_8__23__m2s), .qb(),
		.d(n3468), .sdi(n2596), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__23__slave ( .q(_RegFile_8__23), .qb(n2597), .d(_RegFile_reg_8__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__24__master ( .q(_RegFile_reg_8__24__m2s), .qb(),
		.d(n3469), .sdi(n2597), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__24__slave ( .q(_RegFile_8__24), .qb(n2598), .d(_RegFile_reg_8__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__25__master ( .q(_RegFile_reg_8__25__m2s), .qb(),
		.d(n3470), .sdi(n2598), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__25__slave ( .q(_RegFile_8__25), .qb(n2599), .d(_RegFile_reg_8__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__26__master ( .q(_RegFile_reg_8__26__m2s), .qb(),
		.d(n3471), .sdi(n2599), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__26__slave ( .q(_RegFile_8__26), .qb(n2600), .d(_RegFile_reg_8__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__27__master ( .q(_RegFile_reg_8__27__m2s), .qb(),
		.d(n3472), .sdi(n2600), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__27__slave ( .q(_RegFile_8__27), .qb(n2601), .d(_RegFile_reg_8__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__28__master ( .q(_RegFile_reg_8__28__m2s), .qb(),
		.d(n3473), .sdi(n2601), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n921),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__28__slave ( .q(_RegFile_8__28), .qb(n2602), .d(_RegFile_reg_8__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n921), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__29__master ( .q(_RegFile_reg_8__29__m2s), .qb(),
		.d(n3474), .sdi(n2602), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__29__slave ( .q(_RegFile_8__29), .qb(n2603), .d(_RegFile_reg_8__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__2__master ( .q(_RegFile_reg_8__2__m2s), .qb(),
		.d(n3447), .sdi(n4303), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__2__slave ( .q(_RegFile_8__2), .qb(n4302), .d(_RegFile_reg_8__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__30__master ( .q(_RegFile_reg_8__30__m2s), .qb(),
		.d(n3475), .sdi(n2603), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__30__slave ( .q(_RegFile_8__30), .qb(n2604), .d(_RegFile_reg_8__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__31__master ( .q(_RegFile_reg_8__31__m2s), .qb(),
		.d(n3476), .sdi(n2604), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__31__slave ( .q(_RegFile_8__31), .qb(n2605), .d(_RegFile_reg_8__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__3__master ( .q(_RegFile_reg_8__3__m2s), .qb(),
		.d(n3448), .sdi(n4302), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__3__slave ( .q(_RegFile_8__3), .qb(n4301), .d(_RegFile_reg_8__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__4__master ( .q(_RegFile_reg_8__4__m2s), .qb(),
		.d(n3449), .sdi(n4301), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__4__slave ( .q(_RegFile_8__4), .qb(n4300), .d(_RegFile_reg_8__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__5__master ( .q(_RegFile_reg_8__5__m2s), .qb(),
		.d(n3450), .sdi(n4300), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__5__slave ( .q(_RegFile_8__5), .qb(n4299), .d(_RegFile_reg_8__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__6__master ( .q(_RegFile_reg_8__6__m2s), .qb(),
		.d(n3451), .sdi(n4299), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__6__slave ( .q(_RegFile_8__6), .qb(n4298), .d(_RegFile_reg_8__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__7__master ( .q(_RegFile_reg_8__7__m2s), .qb(),
		.d(n3452), .sdi(n4298), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__7__slave ( .q(_RegFile_8__7), .qb(n4297), .d(_RegFile_reg_8__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__8__master ( .q(_RegFile_reg_8__8__m2s), .qb(),
		.d(n3453), .sdi(n4297), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__8__slave ( .q(_RegFile_8__8), .qb(n2606), .d(_RegFile_reg_8__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_8__9__master ( .q(_RegFile_reg_8__9__m2s), .qb(),
		.d(n3454), .sdi(n2606), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_8__9__slave ( .q(_RegFile_8__9), .qb(n2607), .d(_RegFile_reg_8__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__0__master ( .q(_RegFile_reg_9__0__m2s), .qb(),
		.d(n3413), .sdi(n2605), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__0__slave ( .q(_RegFile_9__0), .qb(n4296), .d(_RegFile_reg_9__0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__10__master ( .q(_RegFile_reg_9__10__m2s), .qb(),
		.d(n3423), .sdi(n2631), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__10__slave ( .q(_RegFile_9__10), .qb(n2608), .d(_RegFile_reg_9__10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__11__master ( .q(_RegFile_reg_9__11__m2s), .qb(),
		.d(n3424), .sdi(n2608), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__11__slave ( .q(_RegFile_9__11), .qb(n2609), .d(_RegFile_reg_9__11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__12__master ( .q(_RegFile_reg_9__12__m2s), .qb(),
		.d(n3425), .sdi(n2609), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n980),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__12__slave ( .q(_RegFile_9__12), .qb(n2610), .d(_RegFile_reg_9__12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n980), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__13__master ( .q(_RegFile_reg_9__13__m2s), .qb(),
		.d(n3426), .sdi(n2610), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__13__slave ( .q(_RegFile_9__13), .qb(n2611), .d(_RegFile_reg_9__13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__14__master ( .q(_RegFile_reg_9__14__m2s), .qb(),
		.d(n3427), .sdi(n2611), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__14__slave ( .q(_RegFile_9__14), .qb(n2612), .d(_RegFile_reg_9__14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__15__master ( .q(_RegFile_reg_9__15__m2s), .qb(),
		.d(n3428), .sdi(n2612), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__15__slave ( .q(_RegFile_9__15), .qb(n2613), .d(_RegFile_reg_9__15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__16__master ( .q(_RegFile_reg_9__16__m2s), .qb(),
		.d(n3429), .sdi(n2613), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__16__slave ( .q(_RegFile_9__16), .qb(n2614), .d(_RegFile_reg_9__16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__17__master ( .q(_RegFile_reg_9__17__m2s), .qb(),
		.d(n3430), .sdi(n2614), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__17__slave ( .q(_RegFile_9__17), .qb(n2615), .d(_RegFile_reg_9__17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__18__master ( .q(_RegFile_reg_9__18__m2s), .qb(),
		.d(n3431), .sdi(n2615), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__18__slave ( .q(_RegFile_9__18), .qb(n2616), .d(_RegFile_reg_9__18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__19__master ( .q(_RegFile_reg_9__19__m2s), .qb(),
		.d(n3432), .sdi(n2616), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__19__slave ( .q(_RegFile_9__19), .qb(n2617), .d(_RegFile_reg_9__19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__1__master ( .q(_RegFile_reg_9__1__m2s), .qb(),
		.d(n3414), .sdi(n4296), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__1__slave ( .q(_RegFile_9__1), .qb(n4295), .d(_RegFile_reg_9__1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__20__master ( .q(_RegFile_reg_9__20__m2s), .qb(),
		.d(n3433), .sdi(n2617), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__20__slave ( .q(_RegFile_9__20), .qb(n2618), .d(_RegFile_reg_9__20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__21__master ( .q(_RegFile_reg_9__21__m2s), .qb(),
		.d(n3434), .sdi(n2618), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__21__slave ( .q(_RegFile_9__21), .qb(n2619), .d(_RegFile_reg_9__21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__22__master ( .q(_RegFile_reg_9__22__m2s), .qb(),
		.d(n3435), .sdi(n2619), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__22__slave ( .q(_RegFile_9__22), .qb(n2620), .d(_RegFile_reg_9__22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__23__master ( .q(_RegFile_reg_9__23__m2s), .qb(),
		.d(n3436), .sdi(n2620), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__23__slave ( .q(_RegFile_9__23), .qb(n2621), .d(_RegFile_reg_9__23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__24__master ( .q(_RegFile_reg_9__24__m2s), .qb(),
		.d(n3437), .sdi(n2621), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__24__slave ( .q(_RegFile_9__24), .qb(n2622), .d(_RegFile_reg_9__24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__25__master ( .q(_RegFile_reg_9__25__m2s), .qb(),
		.d(n3438), .sdi(n2622), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__25__slave ( .q(_RegFile_9__25), .qb(n2623), .d(_RegFile_reg_9__25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__26__master ( .q(_RegFile_reg_9__26__m2s), .qb(),
		.d(n3439), .sdi(n2623), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n920),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__26__slave ( .q(_RegFile_9__26), .qb(n2624), .d(_RegFile_reg_9__26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n920), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__27__master ( .q(_RegFile_reg_9__27__m2s), .qb(),
		.d(n3440), .sdi(n2624), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__27__slave ( .q(_RegFile_9__27), .qb(n2625), .d(_RegFile_reg_9__27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__28__master ( .q(_RegFile_reg_9__28__m2s), .qb(),
		.d(n3441), .sdi(n2625), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__28__slave ( .q(_RegFile_9__28), .qb(n2626), .d(_RegFile_reg_9__28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__29__master ( .q(_RegFile_reg_9__29__m2s), .qb(),
		.d(n3442), .sdi(n2626), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__29__slave ( .q(_RegFile_9__29), .qb(n2627), .d(_RegFile_reg_9__29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__2__master ( .q(_RegFile_reg_9__2__m2s), .qb(),
		.d(n3415), .sdi(n4295), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__2__slave ( .q(_RegFile_9__2), .qb(n4294), .d(_RegFile_reg_9__2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__30__master ( .q(_RegFile_reg_9__30__m2s), .qb(),
		.d(n3443), .sdi(n2627), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__30__slave ( .q(_RegFile_9__30), .qb(n2628), .d(_RegFile_reg_9__30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__31__master ( .q(_RegFile_reg_9__31__m2s), .qb(),
		.d(n3444), .sdi(n2628), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__31__slave ( .q(_RegFile_9__31), .qb(n2629), .d(_RegFile_reg_9__31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__3__master ( .q(_RegFile_reg_9__3__m2s), .qb(),
		.d(n3416), .sdi(n4294), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__3__slave ( .q(_RegFile_9__3), .qb(n4293), .d(_RegFile_reg_9__3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__4__master ( .q(_RegFile_reg_9__4__m2s), .qb(),
		.d(n3417), .sdi(n4293), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__4__slave ( .q(_RegFile_9__4), .qb(n4292), .d(_RegFile_reg_9__4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__5__master ( .q(_RegFile_reg_9__5__m2s), .qb(),
		.d(n3418), .sdi(n4292), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__5__slave ( .q(_RegFile_9__5), .qb(n4291), .d(_RegFile_reg_9__5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__6__master ( .q(_RegFile_reg_9__6__m2s), .qb(),
		.d(n3419), .sdi(n4291), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__6__slave ( .q(_RegFile_9__6), .qb(n4290), .d(_RegFile_reg_9__6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__7__master ( .q(_RegFile_reg_9__7__m2s), .qb(),
		.d(n3420), .sdi(n4290), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__7__slave ( .q(_RegFile_9__7), .qb(n4289), .d(_RegFile_reg_9__7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__8__master ( .q(_RegFile_reg_9__8__m2s), .qb(),
		.d(n3421), .sdi(n4289), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__8__slave ( .q(_RegFile_9__8), .qb(n2630), .d(_RegFile_reg_9__8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 _RegFile_reg_9__9__master ( .q(_RegFile_reg_9__9__m2s), .qb(),
		.d(n3422), .sdi(n2630), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 _RegFile_reg_9__9__slave ( .q(_RegFile_9__9), .qb(n2631), .d(_RegFile_reg_9__9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2), .sync_sel(sync_sel) );
	ID_DW01_sub_32_2_test_1 add_489 ( .A({ NPC[31], NPC[30], NPC[29], NPC[28],
		NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], NPC[21], NPC[20],
		NPC[19], NPC[18], NPC[17], NPC[16], NPC[15], NPC[14], NPC[13], NPC[12],
		NPC[11], NPC[10], NPC[9], NPC[8], NPC[7], NPC[6], NPC[5], NPC[4], NPC[3],
		n737, NPC[1], NPC[0]}), .B({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0,
		1'b0}), .CI(1'b0), .DIFF({ N5350, N5349, N5348, N5347, N5346, N5345,
		N5344, N5343, N5342, N5341, N5340, N5339, N5338, N5337, N5336, N5335,
		N5334, N5333, N5332, N5331, N5330, N5329, N5328, N5327, N5326, N5325,
		N5324, N5323, N5322, N5321, N5320, N5319}), .CO() );
	ID_DW01_sub_32_0_test_1 add_609 ( .A(NPC), .B({ 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .DIFF({ N5418, N5417, N5416, N5415,
		N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406, N5405,
		N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396, N5395,
		N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387}), .CO() );
	ID_DW01_sub_32_1_test_1 add_779 ( .A({ NPC[31], NPC[30], NPC[29], NPC[28],
		NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], NPC[21], NPC[20],
		NPC[19], NPC[18], NPC[17], NPC[16], NPC[15], NPC[14], NPC[13], NPC[12],
		NPC[11], NPC[10], NPC[9], NPC[8], NPC[7], NPC[6], NPC[5], NPC[4], n811,
		n866, NPC[1], NPC[0]}), .B({ 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0,
		1'b0}), .CI(1'b0), .DIFF({ N6017, N6016, N6015, N6014, N6013, N6012,
		N6011, N6010, N6009, N6008, N6007, N6006, N6005, N6004, N6003, N6002,
		N6001, N6000, N5999, N5998, N5997, N5996, N5995, N5994, N5993, N5992,
		N5991, N5990, N5989, N5988, N5987, N5986}), .CO() );
	smlatnr_2 branch_address_reg_0__master ( .q(branch_address_reg_0__m2s),
		.qb(), .d(n3824), .sdi(WB_index_4), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n969), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_0__slave ( .q(branch_address[0]), .qb(n4112),
		.d(branch_address_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_10__master ( .q(branch_address_reg_10__m2s),
		.qb(), .d(n3834), .sdi(n4104), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n969),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_10__slave ( .q(branch_address[10]), .qb(n4103),
		.d(branch_address_reg_10__m2s), .g(Ctrl__Regs_1__en2), .rb(n969), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_11__master ( .q(branch_address_reg_11__m2s),
		.qb(), .d(n3835), .sdi(n4103), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_11__slave ( .q(branch_address[11]), .qb(n4102),
		.d(branch_address_reg_11__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_12__master ( .q(branch_address_reg_12__m2s),
		.qb(), .d(n3836), .sdi(n4102), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_12__slave ( .q(branch_address[12]), .qb(n4101),
		.d(branch_address_reg_12__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_13__master ( .q(branch_address_reg_13__m2s),
		.qb(), .d(n3837), .sdi(n4101), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_13__slave ( .q(branch_address[13]), .qb(n4100),
		.d(branch_address_reg_13__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_14__master ( .q(branch_address_reg_14__m2s),
		.qb(), .d(n3838), .sdi(n4100), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_14__slave ( .q(branch_address[14]), .qb(n4099),
		.d(branch_address_reg_14__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 branch_address_reg_15__master ( .q(branch_address_reg_15__m2s),
		.qb(), .d(n3839), .sdi(n4099), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 branch_address_reg_15__slave ( .q(branch_address[15]), .qb(n4098),
		.d(branch_address_reg_15__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_16__master ( .q(branch_address_reg_16__m2s),
		.qb(), .d(n3840), .sdi(n4098), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_16__slave ( .q(branch_address[16]), .qb(n4097),
		.d(branch_address_reg_16__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_17__master ( .q(branch_address_reg_17__m2s),
		.qb(), .d(n3841), .sdi(n4097), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_17__slave ( .q(branch_address[17]), .qb(n4096),
		.d(branch_address_reg_17__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_18__master ( .q(branch_address_reg_18__m2s),
		.qb(), .d(n3842), .sdi(n4096), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_18__slave ( .q(branch_address[18]), .qb(n4095),
		.d(branch_address_reg_18__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_19__master ( .q(branch_address_reg_19__m2s),
		.qb(), .d(n3843), .sdi(n4095), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_19__slave ( .q(branch_address[19]), .qb(n4094),
		.d(branch_address_reg_19__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 branch_address_reg_1__master ( .q(branch_address_reg_1__m2s),
		.qb(), .d(n3825), .sdi(n4112), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 branch_address_reg_1__slave ( .q(branch_address[1]), .qb(n4111),
		.d(branch_address_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_20__master ( .q(branch_address_reg_20__m2s),
		.qb(), .d(n3844), .sdi(n4094), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_20__slave ( .q(branch_address[20]), .qb(n4093),
		.d(branch_address_reg_20__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_21__master ( .q(branch_address_reg_21__m2s),
		.qb(), .d(n3845), .sdi(n4093), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_21__slave ( .q(branch_address[21]), .qb(n4092),
		.d(branch_address_reg_21__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_22__master ( .q(branch_address_reg_22__m2s),
		.qb(), .d(n3846), .sdi(n4092), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_22__slave ( .q(branch_address[22]), .qb(n4091),
		.d(branch_address_reg_22__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_23__master ( .q(branch_address_reg_23__m2s),
		.qb(), .d(n3847), .sdi(n4091), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_23__slave ( .q(branch_address[23]), .qb(n4090),
		.d(branch_address_reg_23__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_24__master ( .q(branch_address_reg_24__m2s),
		.qb(), .d(n3848), .sdi(n4090), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n919),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_24__slave ( .q(branch_address[24]), .qb(n4089),
		.d(branch_address_reg_24__m2s), .g(Ctrl__Regs_1__en2), .rb(n919), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_25__master ( .q(branch_address_reg_25__m2s),
		.qb(), .d(n3849), .sdi(n4089), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_25__slave ( .q(branch_address[25]), .qb(n4088),
		.d(branch_address_reg_25__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_26__master ( .q(branch_address_reg_26__m2s),
		.qb(), .d(n3850), .sdi(n4088), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_26__slave ( .q(branch_address[26]), .qb(n4087),
		.d(branch_address_reg_26__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 branch_address_reg_27__master ( .q(branch_address_reg_27__m2s),
		.qb(), .d(n3851), .sdi(n4087), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 branch_address_reg_27__slave ( .q(branch_address[27]), .qb(n4086),
		.d(branch_address_reg_27__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_28__master ( .q(branch_address_reg_28__m2s),
		.qb(), .d(n3852), .sdi(n4086), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_28__slave ( .q(branch_address[28]), .qb(n4085),
		.d(branch_address_reg_28__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_29__master ( .q(branch_address_reg_29__m2s),
		.qb(), .d(n3853), .sdi(n4085), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_29__slave ( .q(branch_address[29]), .qb(n4084),
		.d(branch_address_reg_29__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_2__master ( .q(branch_address_reg_2__m2s),
		.qb(), .d(n3826), .sdi(n4111), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_2__slave ( .q(branch_address[2]), .qb(n4110),
		.d(branch_address_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_30__master ( .q(branch_address_reg_30__m2s),
		.qb(), .d(n3854), .sdi(n4084), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_30__slave ( .q(branch_address[30]), .qb(n4083),
		.d(branch_address_reg_30__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_31__master ( .q(branch_address_reg_31__m2s),
		.qb(), .d(_branch_address_reg_31_net46811), .sdi(n4083), .se(test_se),
		.g(Ctrl__Regs_1__en1), .rb(n918), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_31__slave ( .q(branch_address[31]), .qb(n2632),
		.d(branch_address_reg_31__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_3__master ( .q(branch_address_reg_3__m2s),
		.qb(), .d(n3827), .sdi(n4110), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_3__slave ( .q(branch_address[3]), .qb(n4109),
		.d(branch_address_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_4__master ( .q(branch_address_reg_4__m2s),
		.qb(), .d(n3828), .sdi(n4109), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_4__slave ( .q(branch_address[4]), .qb(n4108),
		.d(branch_address_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_5__master ( .q(branch_address_reg_5__m2s),
		.qb(), .d(n3829), .sdi(n4108), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_5__slave ( .q(branch_address[5]), .qb(n4107),
		.d(branch_address_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_6__master ( .q(branch_address_reg_6__m2s),
		.qb(), .d(n3830), .sdi(n4107), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n981),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_6__slave ( .q(branch_address[6]), .qb(n4106),
		.d(branch_address_reg_6__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_7__master ( .q(branch_address_reg_7__m2s),
		.qb(), .d(n3831), .sdi(n4106), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_7__slave ( .q(branch_address[7]), .qb(n2633),
		.d(branch_address_reg_7__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_8__master ( .q(branch_address_reg_8__m2s),
		.qb(), .d(n3832), .sdi(branch_address[7]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n981), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_8__slave ( .q(branch_address[8]), .qb(n4105),
		.d(branch_address_reg_8__m2s), .g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_address_reg_9__master ( .q(branch_address_reg_9__m2s),
		.qb(), .d(n3833), .sdi(n4105), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_address_reg_9__slave ( .q(branch_address[9]), .qb(n4104),
		.d(branch_address_reg_9__m2s), .g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_2 branch_sig_reg__master ( .q(branch_sig_reg__m2s), .qb(), .d(n3823),
		.sdi(branch_address[31]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 branch_sig_reg__slave ( .q(branch_sig), .qb(n2634), .d(branch_sig_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 counter_reg_0__master ( .q(counter_reg_0__m2s), .qb(), .d(_counter_reg_0_net48671),
		.sdi(n2634), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 counter_reg_0__slave ( .q(n3950), .qb(n787), .d(counter_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 counter_reg_1__master ( .q(counter_reg_1__m2s), .qb(), .d(_counter_reg_1_net48651),
		.sdi(counter[0]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 counter_reg_1__slave ( .q(n3949), .qb(n780), .d(counter_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_0__master ( .q(current_IR_reg_0__m2s), .qb(),
		.d(n3733), .sdi(n790), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_0__slave ( .q(current_IR_0), .qb(n4082), .d(current_IR_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_10__master ( .q(current_IR_reg_10__m2s), .qb(),
		.d(n3742), .sdi(n629), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_10__slave ( .q(current_IR_10), .qb(n632), .d(current_IR_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_11__master ( .q(current_IR_reg_11__m2s), .qb(),
		.d(n3743), .sdi(n632), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_11__slave ( .q(n4076), .qb(n571), .d(current_IR_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_12__master ( .q(current_IR_reg_12__m2s), .qb(),
		.d(n3744), .sdi(n4076), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_12__slave ( .q(n4075), .qb(n652), .d(current_IR_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_13__master ( .q(current_IR_reg_13__m2s), .qb(),
		.d(n3745), .sdi(n4075), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_13__slave ( .q(n4074), .qb(n570), .d(current_IR_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_14__master ( .q(current_IR_reg_14__m2s), .qb(),
		.d(n3746), .sdi(n4074), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_14__slave ( .q(n4073), .qb(n569), .d(current_IR_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_15__master ( .q(current_IR_reg_15__m2s), .qb(),
		.d(n3747), .sdi(n4073), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_15__slave ( .q(n4072), .qb(n568), .d(current_IR_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_16__master ( .q(current_IR_reg_16__m2s), .qb(),
		.d(n3748), .sdi(n4072), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_16__slave ( .q(n644), .qb(n645), .d(current_IR_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_17__master ( .q(current_IR_reg_17__m2s), .qb(),
		.d(n3749), .sdi(n645), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_17__slave ( .q(current_IR_17), .qb(n4071), .d(current_IR_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_18__master ( .q(current_IR_reg_18__m2s), .qb(),
		.d(n3750), .sdi(n4071), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_18__slave ( .q(current_IR_18), .qb(n4070), .d(current_IR_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_19__master ( .q(current_IR_reg_19__m2s), .qb(),
		.d(n3751), .sdi(n4070), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_19__slave ( .q(current_IR_19), .qb(n657), .d(current_IR_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_1__master ( .q(current_IR_reg_1__m2s), .qb(),
		.d(_current_IR_reg_1_net49291), .sdi(n4082), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n981), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_1__slave ( .q(current_IR_1), .qb(n4081), .d(current_IR_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n981), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_20__master ( .q(current_IR_reg_20__m2s), .qb(),
		.d(n3752), .sdi(n657), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_20__slave ( .q(n4069), .qb(n567), .d(current_IR_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_21__master ( .q(current_IR_reg_21__m2s), .qb(),
		.d(n3753), .sdi(n4069), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_21__slave ( .q(current_IR_21), .qb(n646), .d(current_IR_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_22__master ( .q(current_IR_reg_22__m2s), .qb(),
		.d(n3754), .sdi(n646), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_22__slave ( .q(n660), .qb(n661), .d(current_IR_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_23__master ( .q(current_IR_reg_23__m2s), .qb(),
		.d(n3755), .sdi(n661), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_23__slave ( .q(current_IR_23), .qb(n659), .d(current_IR_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_24__master ( .q(current_IR_reg_24__m2s), .qb(),
		.d(n3756), .sdi(n659), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_24__slave ( .q(current_IR_24), .qb(n4068), .d(current_IR_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_25__master ( .q(current_IR_reg_25__m2s), .qb(),
		.d(n3757), .sdi(n4068), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_25__slave ( .q(n4067), .qb(n666), .d(current_IR_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_26__master ( .q(current_IR_reg_26__m2s), .qb(),
		.d(n3758), .sdi(n4067), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_26__slave ( .q(n4066), .qb(n852), .d(current_IR_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_27__master ( .q(current_IR_reg_27__m2s), .qb(),
		.d(n3759), .sdi(n4066), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_27__slave ( .q(current_IR_27), .qb(n4065), .d(current_IR_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_28__master ( .q(current_IR_reg_28__m2s), .qb(),
		.d(n3760), .sdi(n4065), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_28__slave ( .q(n4064), .qb(n566), .d(current_IR_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_29__master ( .q(current_IR_reg_29__m2s), .qb(),
		.d(n3761), .sdi(n4064), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_29__slave ( .q(current_IR_29), .qb(n656), .d(current_IR_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_2__master ( .q(current_IR_reg_2__m2s), .qb(),
		.d(n3734), .sdi(n4081), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n918),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_2__slave ( .q(current_IR_2), .qb(n4080), .d(current_IR_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n918), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_30__master ( .q(current_IR_reg_30__m2s), .qb(),
		.d(n3762), .sdi(n656), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_30__slave ( .q(current_IR_30), .qb(n658), .d(current_IR_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_31__master ( .q(current_IR_reg_31__m2s), .qb(),
		.d(n3763), .sdi(n658), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_31__slave ( .q(current_IR_31), .qb(n633), .d(current_IR_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_3__master ( .q(current_IR_reg_3__m2s), .qb(),
		.d(n3735), .sdi(n4080), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n948),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_3__slave ( .q(current_IR_3), .qb(n651), .d(current_IR_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n948), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_4__master ( .q(current_IR_reg_4__m2s), .qb(),
		.d(n3736), .sdi(n651), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_4__slave ( .q(current_IR_4), .qb(n4079), .d(current_IR_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_5__master ( .q(current_IR_reg_5__m2s), .qb(),
		.d(n3737), .sdi(n4079), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_5__slave ( .q(n4078), .qb(n565), .d(current_IR_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_6__master ( .q(current_IR_reg_6__m2s), .qb(),
		.d(n3738), .sdi(n4078), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_6__slave ( .q(current_IR_6), .qb(n631), .d(current_IR_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_7__master ( .q(current_IR_reg_7__m2s), .qb(),
		.d(n3739), .sdi(n631), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_7__slave ( .q(current_IR_7), .qb(n4077), .d(current_IR_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_8__master ( .q(current_IR_reg_8__m2s), .qb(),
		.d(n3740), .sdi(n4077), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_8__slave ( .q(current_IR_8), .qb(n630), .d(current_IR_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 current_IR_reg_9__master ( .q(current_IR_reg_9__m2s), .qb(),
		.d(n3741), .sdi(n630), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n938),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 current_IR_reg_9__slave ( .q(current_IR_9), .qb(n629), .d(current_IR_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n938), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 delay_slot_reg__master ( .q(delay_slot_reg__m2s), .qb(), .d(n2707),
		.sdi(n633), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 delay_slot_reg__slave ( .q(delay_slot), .qb(n883), .d(delay_slot_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 intr_slot_reg__master ( .q(intr_slot_reg__m2s), .qb(), .d(n2640),
		.sdi(n883), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 intr_slot_reg__slave ( .q(intr_slot), .qb(n564), .d(intr_slot_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 mem_read_reg__master ( .q(mem_read_reg__m2s), .qb(), .d(n3777),
		.sdi(intr_slot), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 mem_read_reg__slave ( .q(mem_read), .qb(n2635), .d(mem_read_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 mem_to_reg_reg__master ( .q(mem_to_reg_reg__m2s), .qb(), .d(n3778),
		.sdi(mem_read), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 mem_to_reg_reg__slave ( .q(mem_to_reg), .qb(n2636), .d(mem_to_reg_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 mem_write_reg__master ( .q(mem_write_reg__m2s), .qb(), .d(n3776),
		.sdi(mem_to_reg), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 mem_write_reg__slave ( .q(mem_write), .qb(n2637), .d(mem_write_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 opcode_of_MEM_reg_0__master ( .q(opcode_of_MEM_reg_0__m2s), .qb(),
		.d(IR_opcode_field[0]), .sdi(mem_write), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_MEM_reg_0__slave ( .q(opcode_of_MEM_0), .qb(n3924),
		.d(opcode_of_MEM_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 opcode_of_MEM_reg_1__master ( .q(opcode_of_MEM_reg_1__m2s), .qb(),
		.d(IR_opcode_field[1]), .sdi(opcode_of_MEM_0), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_MEM_reg_1__slave ( .q(opcode_of_MEM_1), .qb(n4063),
		.d(opcode_of_MEM_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 opcode_of_MEM_reg_2__master ( .q(opcode_of_MEM_reg_2__m2s), .qb(),
		.d(IR_opcode_field[2]), .sdi(n4063), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_MEM_reg_2__slave ( .q(opcode_of_MEM_2), .qb(n3933),
		.d(opcode_of_MEM_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 opcode_of_MEM_reg_3__master ( .q(opcode_of_MEM_reg_3__m2s), .qb(),
		.d(IR_opcode_field[3]), .sdi(n3933), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_MEM_reg_3__slave ( .q(opcode_of_MEM_3), .qb(n3932),
		.d(opcode_of_MEM_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 opcode_of_MEM_reg_4__master ( .q(opcode_of_MEM_reg_4__m2s), .qb(),
		.d(IR_opcode_field[4]), .sdi(opcode_of_MEM_3), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n911), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 opcode_of_MEM_reg_4__slave ( .q(opcode_of_MEM_4), .qb(n4062),
		.d(opcode_of_MEM_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 opcode_of_MEM_reg_5__master ( .q(opcode_of_MEM_reg_5__m2s), .qb(),
		.d(IR_opcode_field[5]), .sdi(n4062), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_MEM_reg_5__slave ( .q(opcode_of_MEM_5), .qb(n4061),
		.d(opcode_of_MEM_reg_5__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 opcode_of_WB_reg_0__master ( .q(opcode_of_WB_reg_0__m2s), .qb(),
		.d(opcode_of_MEM_0), .sdi(n4061), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_WB_reg_0__slave ( .q(N13832), .qb(n4060), .d(opcode_of_WB_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 opcode_of_WB_reg_1__master ( .q(opcode_of_WB_reg_1__m2s), .qb(),
		.d(opcode_of_MEM_1), .sdi(n4060), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_WB_reg_1__slave ( .q(n4059), .qb(n3887), .d(opcode_of_WB_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 opcode_of_WB_reg_2__master ( .q(opcode_of_WB_reg_2__m2s), .qb(),
		.d(opcode_of_MEM_2), .sdi(n4059), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_WB_reg_2__slave ( .q(n3888), .qb(n4058), .d(opcode_of_WB_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 opcode_of_WB_reg_3__master ( .q(opcode_of_WB_reg_3__m2s), .qb(),
		.d(opcode_of_MEM_3), .sdi(n4058), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_WB_reg_3__slave ( .q(n4057), .qb(n3889), .d(opcode_of_WB_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 opcode_of_WB_reg_4__master ( .q(opcode_of_WB_reg_4__m2s), .qb(),
		.d(opcode_of_MEM_4), .sdi(n4057), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n912), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_WB_reg_4__slave ( .q(n4056), .qb(n3890), .d(opcode_of_WB_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 opcode_of_WB_reg_5__master ( .q(opcode_of_WB_reg_5__m2s), .qb(),
		.d(opcode_of_MEM_5), .sdi(n4056), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 opcode_of_WB_reg_5__slave ( .q(opcode_of_WB_5), .qb(n4055), .d(opcode_of_WB_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rd_addr_reg_0__master ( .q(rd_addr_reg_0__m2s), .qb(), .d(n3781),
		.sdi(n4055), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rd_addr_reg_0__slave ( .q(rd_addr[0]), .qb(n669), .d(rd_addr_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rd_addr_reg_1__master ( .q(rd_addr_reg_1__m2s), .qb(), .d(n3782),
		.sdi(rd_addr[0]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rd_addr_reg_1__slave ( .q(rd_addr[1]), .qb(n563), .d(rd_addr_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rd_addr_reg_2__master ( .q(rd_addr_reg_2__m2s), .qb(), .d(n3783),
		.sdi(rd_addr[1]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rd_addr_reg_2__slave ( .q(rd_addr[2]), .qb(n670), .d(rd_addr_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rd_addr_reg_3__master ( .q(rd_addr_reg_3__m2s), .qb(), .d(n3784),
		.sdi(rd_addr[2]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rd_addr_reg_3__slave ( .q(rd_addr[3]), .qb(n4054), .d(rd_addr_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rd_addr_reg_4__master ( .q(rd_addr_reg_4__m2s), .qb(), .d(n3785),
		.sdi(n4054), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rd_addr_reg_4__slave ( .q(rd_addr[4]), .qb(n562), .d(rd_addr_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_dst_of_MEM_reg_0__master ( .q(reg_dst_of_MEM_reg_0__m2s),
		.qb(), .d(reg_dst_of_EX_0), .sdi(rd_addr[4]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_dst_of_MEM_reg_0__slave ( .q(reg_dst_of_MEM_0), .qb(n4053),
		.d(reg_dst_of_MEM_reg_0__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_dst_of_MEM_reg_1__master ( .q(reg_dst_of_MEM_reg_1__m2s),
		.qb(), .d(reg_dst_of_EX_1), .sdi(n4053), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_1 reg_dst_of_MEM_reg_1__slave ( .q(reg_dst_of_MEM_1), .qb(n4052),
		.d(reg_dst_of_MEM_reg_1__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_dst_of_MEM_reg_2__master ( .q(reg_dst_of_MEM_reg_2__m2s),
		.qb(), .d(reg_dst_of_EX_2), .sdi(n4052), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n913), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_dst_of_MEM_reg_2__slave ( .q(reg_dst_of_MEM_2), .qb(n655),
		.d(reg_dst_of_MEM_reg_2__m2s), .g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_dst_of_MEM_reg_3__master ( .q(reg_dst_of_MEM_reg_3__m2s),
		.qb(), .d(reg_dst_of_EX_3), .sdi(reg_dst_of_MEM_2), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_dst_of_MEM_reg_3__slave ( .q(reg_dst_of_MEM_3), .qb(n634),
		.d(reg_dst_of_MEM_reg_3__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_dst_of_MEM_reg_4__master ( .q(reg_dst_of_MEM_reg_4__m2s),
		.qb(), .d(reg_dst_of_EX_4), .sdi(reg_dst_of_MEM_3), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n914), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_dst_of_MEM_reg_4__slave ( .q(reg_dst_of_MEM_4), .qb(n635),
		.d(reg_dst_of_MEM_reg_4__m2s), .g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2),
		.sync_sel(sync_sel) );
	smlatnr_1 reg_dst_reg__master ( .q(reg_dst_reg__m2s), .qb(), .d(n3780),
		.sdi(reg_dst_of_MEM_4), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_dst_reg__slave ( .q(reg_dst), .qb(n703), .d(reg_dst_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_0__master ( .q(reg_out_A_reg_0__m2s), .qb(), .d(N6718),
		.sdi(n703), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_0__slave ( .q(reg_out_A[0]), .qb(n4051), .d(reg_out_A_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_10__master ( .q(reg_out_A_reg_10__m2s), .qb(),
		.d(N6728), .sdi(n4042), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_10__slave ( .q(n3968), .qb(n4041), .d(reg_out_A_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_11__master ( .q(reg_out_A_reg_11__m2s), .qb(),
		.d(N6729), .sdi(n4041), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_11__slave ( .q(n3967), .qb(n4040), .d(reg_out_A_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_12__master ( .q(reg_out_A_reg_12__m2s), .qb(),
		.d(N6730), .sdi(n4040), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_12__slave ( .q(n3966), .qb(n4039), .d(reg_out_A_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_13__master ( .q(reg_out_A_reg_13__m2s), .qb(),
		.d(N6731), .sdi(n4039), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_13__slave ( .q(reg_out_A[13]), .qb(n4038), .d(reg_out_A_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_14__master ( .q(reg_out_A_reg_14__m2s), .qb(),
		.d(N6732), .sdi(n4038), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_14__slave ( .q(reg_out_A[14]), .qb(n4037), .d(reg_out_A_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_15__master ( .q(reg_out_A_reg_15__m2s), .qb(),
		.d(N6733), .sdi(n4037), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_15__slave ( .q(reg_out_A[15]), .qb(n4036), .d(reg_out_A_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_16__master ( .q(reg_out_A_reg_16__m2s), .qb(),
		.d(N6734), .sdi(n4036), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_16__slave ( .q(n3965), .qb(n4035), .d(reg_out_A_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_17__master ( .q(reg_out_A_reg_17__m2s), .qb(),
		.d(N6735), .sdi(n4035), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_17__slave ( .q(n3964), .qb(n4034), .d(reg_out_A_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_18__master ( .q(reg_out_A_reg_18__m2s), .qb(),
		.d(N6736), .sdi(n4034), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_18__slave ( .q(n3963), .qb(n4033), .d(reg_out_A_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_19__master ( .q(reg_out_A_reg_19__m2s), .qb(),
		.d(N6737), .sdi(n4033), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_19__slave ( .q(n3962), .qb(n4032), .d(reg_out_A_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_1__master ( .q(reg_out_A_reg_1__m2s), .qb(), .d(N6719),
		.sdi(n4051), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_1__slave ( .q(reg_out_A[1]), .qb(n4050), .d(reg_out_A_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_20__master ( .q(reg_out_A_reg_20__m2s), .qb(),
		.d(N6738), .sdi(n4032), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_20__slave ( .q(n3961), .qb(n4031), .d(reg_out_A_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_21__master ( .q(reg_out_A_reg_21__m2s), .qb(),
		.d(N6739), .sdi(n4031), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_21__slave ( .q(n3960), .qb(n4030), .d(reg_out_A_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_22__master ( .q(reg_out_A_reg_22__m2s), .qb(),
		.d(N6740), .sdi(n4030), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_22__slave ( .q(n3959), .qb(n4029), .d(reg_out_A_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_23__master ( .q(reg_out_A_reg_23__m2s), .qb(),
		.d(N6741), .sdi(n4029), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_23__slave ( .q(n3958), .qb(n4028), .d(reg_out_A_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_24__master ( .q(reg_out_A_reg_24__m2s), .qb(),
		.d(N6742), .sdi(n4028), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n913),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_24__slave ( .q(n3957), .qb(n4027), .d(reg_out_A_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n913), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_25__master ( .q(reg_out_A_reg_25__m2s), .qb(),
		.d(N6743), .sdi(n4027), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_25__slave ( .q(n3956), .qb(n4026), .d(reg_out_A_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_26__master ( .q(reg_out_A_reg_26__m2s), .qb(),
		.d(N6744), .sdi(n4026), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n914),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_26__slave ( .q(n3955), .qb(n4025), .d(reg_out_A_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n914), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_27__master ( .q(reg_out_A_reg_27__m2s), .qb(),
		.d(N6745), .sdi(n4025), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_27__slave ( .q(n3954), .qb(n4024), .d(reg_out_A_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_28__master ( .q(reg_out_A_reg_28__m2s), .qb(),
		.d(N6746), .sdi(n4024), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_28__slave ( .q(n3953), .qb(n4023), .d(reg_out_A_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_29__master ( .q(reg_out_A_reg_29__m2s), .qb(),
		.d(N6747), .sdi(n4023), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_29__slave ( .q(n3952), .qb(n4022), .d(reg_out_A_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_2__master ( .q(reg_out_A_reg_2__m2s), .qb(), .d(N6720),
		.sdi(n4050), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_2__slave ( .q(reg_out_A[2]), .qb(n4049), .d(reg_out_A_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_30__master ( .q(reg_out_A_reg_30__m2s), .qb(),
		.d(N6748), .sdi(n4022), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_30__slave ( .q(n3951), .qb(n4021), .d(reg_out_A_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_A_reg_31__master ( .q(reg_out_A_reg_31__m2s), .qb(),
		.d(N6749), .sdi(n4021), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_A_reg_31__slave ( .q(reg_out_A[31]), .qb(n4020), .d(reg_out_A_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_3__master ( .q(reg_out_A_reg_3__m2s), .qb(), .d(N6721),
		.sdi(n4049), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_3__slave ( .q(n3974), .qb(n4048), .d(reg_out_A_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_4__master ( .q(reg_out_A_reg_4__m2s), .qb(), .d(N6722),
		.sdi(n4048), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_4__slave ( .q(n3973), .qb(n4047), .d(reg_out_A_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_5__master ( .q(reg_out_A_reg_5__m2s), .qb(), .d(N6723),
		.sdi(n4047), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_5__slave ( .q(n3972), .qb(n4046), .d(reg_out_A_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_6__master ( .q(reg_out_A_reg_6__m2s), .qb(), .d(N6724),
		.sdi(n4046), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_6__slave ( .q(reg_out_A[6]), .qb(n4045), .d(reg_out_A_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_7__master ( .q(reg_out_A_reg_7__m2s), .qb(), .d(N6725),
		.sdi(n4045), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_7__slave ( .q(n3971), .qb(n4044), .d(reg_out_A_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_8__master ( .q(reg_out_A_reg_8__m2s), .qb(), .d(N6726),
		.sdi(n4044), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n949), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_A_reg_8__slave ( .q(n3970), .qb(n4043), .d(reg_out_A_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n949), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_A_reg_9__master ( .q(reg_out_A_reg_9__m2s), .qb(), .d(N6727),
		.sdi(n4043), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n915), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 reg_out_A_reg_9__slave ( .q(n3969), .qb(n4042), .d(reg_out_A_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n915), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_0__master ( .q(reg_out_B_reg_0__m2s), .qb(), .d(n4392),
		.sdi(n4020), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_0__slave ( .q(n4458), .qb(n4393), .d(reg_out_B_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_10__master ( .q(reg_out_B_reg_10__m2s), .qb(),
		.d(n4412), .sdi(n4389), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_10__slave ( .q(reg_out_B[10]), .qb(n4413), .d(reg_out_B_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_11__master ( .q(reg_out_B_reg_11__m2s), .qb(),
		.d(n4394), .sdi(n4413), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_11__slave ( .q(reg_out_B[11]), .qb(n4395), .d(reg_out_B_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_12__master ( .q(reg_out_B_reg_12__m2s), .qb(),
		.d(n4432), .sdi(n4395), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_12__slave ( .q(n3979), .qb(n4433), .d(reg_out_B_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_13__master ( .q(reg_out_B_reg_13__m2s), .qb(),
		.d(n4424), .sdi(n4433), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_13__slave ( .q(reg_out_B[13]), .qb(n4425), .d(reg_out_B_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_14__master ( .q(reg_out_B_reg_14__m2s), .qb(),
		.d(n4420), .sdi(n4425), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_14__slave ( .q(reg_out_B[14]), .qb(n4421), .d(reg_out_B_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_15__master ( .q(reg_out_B_reg_15__m2s), .qb(),
		.d(n4402), .sdi(n4421), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_15__slave ( .q(reg_out_B[15]), .qb(n4403), .d(reg_out_B_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_16__master ( .q(reg_out_B_reg_16__m2s), .qb(),
		.d(n4410), .sdi(n4403), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_16__slave ( .q(reg_out_B[16]), .qb(n4411), .d(reg_out_B_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_17__master ( .q(reg_out_B_reg_17__m2s), .qb(),
		.d(n4442), .sdi(n4411), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_17__slave ( .q(n3978), .qb(n4443), .d(reg_out_B_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_18__master ( .q(reg_out_B_reg_18__m2s), .qb(),
		.d(n4426), .sdi(n4443), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_18__slave ( .q(reg_out_B[18]), .qb(n4427), .d(reg_out_B_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_19__master ( .q(reg_out_B_reg_19__m2s), .qb(),
		.d(n4422), .sdi(n4427), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_19__slave ( .q(n4456), .qb(n4423), .d(reg_out_B_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_1__master ( .q(reg_out_B_reg_1__m2s), .qb(), .d(n4444),
		.sdi(n4393), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_reg_1__slave ( .q(n3983), .qb(n4445), .d(reg_out_B_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_20__master ( .q(reg_out_B_reg_20__m2s), .qb(),
		.d(n4390), .sdi(n4423), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_20__slave ( .q(reg_out_B[20]), .qb(n4391), .d(reg_out_B_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_21__master ( .q(reg_out_B_reg_21__m2s), .qb(),
		.d(n4436), .sdi(n4391), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_21__slave ( .q(reg_out_B[21]), .qb(n4437), .d(reg_out_B_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_22__master ( .q(reg_out_B_reg_22__m2s), .qb(),
		.d(n4446), .sdi(n4437), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_22__slave ( .q(n3977), .qb(n4447), .d(reg_out_B_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_23__master ( .q(reg_out_B_reg_23__m2s), .qb(),
		.d(n4414), .sdi(n4447), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_23__slave ( .q(reg_out_B[23]), .qb(n4415), .d(reg_out_B_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_24__master ( .q(reg_out_B_reg_24__m2s), .qb(),
		.d(n4416), .sdi(n4415), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_24__slave ( .q(reg_out_B[24]), .qb(n4417), .d(reg_out_B_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_25__master ( .q(reg_out_B_reg_25__m2s), .qb(),
		.d(n4434), .sdi(n4417), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_25__slave ( .q(n4455), .qb(n4435), .d(reg_out_B_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_26__master ( .q(reg_out_B_reg_26__m2s), .qb(),
		.d(n4406), .sdi(n4435), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_26__slave ( .q(reg_out_B[26]), .qb(n4407), .d(reg_out_B_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_27__master ( .q(reg_out_B_reg_27__m2s), .qb(),
		.d(n4430), .sdi(n4407), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_27__slave ( .q(reg_out_B[27]), .qb(n4431), .d(reg_out_B_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_28__master ( .q(reg_out_B_reg_28__m2s), .qb(),
		.d(n4400), .sdi(n4431), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_28__slave ( .q(reg_out_B[28]), .qb(n4401), .d(reg_out_B_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_29__master ( .q(reg_out_B_reg_29__m2s), .qb(),
		.d(n4396), .sdi(n4401), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n910),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_29__slave ( .q(reg_out_B[29]), .qb(n4397), .d(reg_out_B_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n910), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_2__master ( .q(reg_out_B_reg_2__m2s), .qb(), .d(n4438),
		.sdi(n4445), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_2__slave ( .q(n3982), .qb(n4439), .d(reg_out_B_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_30__master ( .q(reg_out_B_reg_30__m2s), .qb(),
		.d(n4448), .sdi(n4397), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_30__slave ( .q(reg_out_B[30]), .qb(n4449), .d(reg_out_B_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_31__master ( .q(reg_out_B_reg_31__m2s), .qb(),
		.d(n4450), .sdi(n4449), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n911),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_31__slave ( .q(reg_out_B[31]), .qb(n4451), .d(reg_out_B_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n911), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_3__master ( .q(reg_out_B_reg_3__m2s), .qb(), .d(n4440),
		.sdi(n4439), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_reg_3__slave ( .q(n3981), .qb(n4441), .d(reg_out_B_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_4__master ( .q(reg_out_B_reg_4__m2s), .qb(), .d(n4398),
		.sdi(n4441), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n912), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 reg_out_B_reg_4__slave ( .q(n3980), .qb(n4399), .d(reg_out_B_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n912), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_5__master ( .q(reg_out_B_reg_5__m2s), .qb(), .d(n4418),
		.sdi(n4399), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_5__slave ( .q(reg_out_B[5]), .qb(n4419), .d(reg_out_B_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_6__master ( .q(reg_out_B_reg_6__m2s), .qb(), .d(n4404),
		.sdi(n4419), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_reg_6__slave ( .q(n4457), .qb(n4405), .d(reg_out_B_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_reg_7__master ( .q(reg_out_B_reg_7__m2s), .qb(), .d(n4428),
		.sdi(n4405), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 reg_out_B_reg_7__slave ( .q(reg_out_B[7]), .qb(n4429), .d(reg_out_B_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_8__master ( .q(reg_out_B_reg_8__m2s), .qb(), .d(n4408),
		.sdi(n4429), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_8__slave ( .q(reg_out_B[8]), .qb(n4409), .d(reg_out_B_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 reg_out_B_reg_9__master ( .q(reg_out_B_reg_9__m2s), .qb(), .d(n4388),
		.sdi(n4409), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n909), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_8 reg_out_B_reg_9__slave ( .q(reg_out_B[9]), .qb(n4389), .d(reg_out_B_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n909), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_write_reg__master ( .q(reg_write_reg__m2s), .qb(), .d(n3779),
		.sdi(n4451), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 reg_write_reg__slave ( .q(reg_write), .qb(n2638), .d(reg_write_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rt_addr_reg_0__master ( .q(rt_addr_reg_0__m2s), .qb(), .d(n3786),
		.sdi(reg_write), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rt_addr_reg_0__slave ( .q(rt_addr[0]), .qb(n561), .d(rt_addr_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rt_addr_reg_1__master ( .q(rt_addr_reg_1__m2s), .qb(), .d(n3787),
		.sdi(rt_addr[0]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rt_addr_reg_1__slave ( .q(rt_addr[1]), .qb(n560), .d(rt_addr_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rt_addr_reg_2__master ( .q(rt_addr_reg_2__m2s), .qb(), .d(n3788),
		.sdi(rt_addr[1]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n917), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rt_addr_reg_2__slave ( .q(rt_addr[2]), .qb(n559), .d(rt_addr_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n917), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rt_addr_reg_3__master ( .q(rt_addr_reg_3__m2s), .qb(), .d(n3789),
		.sdi(rt_addr[2]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rt_addr_reg_3__slave ( .q(rt_addr[3]), .qb(n671), .d(rt_addr_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 rt_addr_reg_4__master ( .q(rt_addr_reg_4__m2s), .qb(), .d(n3790),
		.sdi(n671), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 rt_addr_reg_4__slave ( .q(rt_addr[4]), .qb(n558), .d(rt_addr_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 slot_num_reg_0__master ( .q(slot_num_reg_0__m2s), .qb(), .d(n2705),
		.sdi(rt_addr[4]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 slot_num_reg_0__slave ( .q(slot_num_0), .qb(n4019), .d(slot_num_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 slot_num_reg_1__master ( .q(slot_num_reg_1__m2s), .qb(), .d(n2706),
		.sdi(n4019), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n916), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 slot_num_reg_1__slave ( .q(slot_num_1), .qb(n557), .d(slot_num_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n916), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 stall_reg__master ( .q(stall_reg__m2s), .qb(), .d(n2708), .sdi(n557),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n982), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 stall_reg__slave ( .q(test_so), .qb(n2639), .d(stall_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n982), .glob_g(global_g2), .sync_sel(sync_sel) );
	ID_DW01_add_32_0_test_1 sub_489 ( .A({ n331, n331, n331, n331, n331, n331,
		n331, n824, n695, n3990, n3998, n802, n337, n878, n892, n340, n887, IR_latched_14,
		IR_latched_13, IR_latched_12, IR_latched_11, IR_latched_10, n809, IR_latched_8,
		n817, n3999, n888, n832, IR_latched_3, IR_latched_2, IR_latched_1, IR_latched_0}),
		.B({ N5350, N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341,
		N5340, N5339, N5338, N5337, N5336, N5335, N5334, N5333, N5332, N5331,
		N5330, N5329, N5328, N5327, N5326, N5325, N5324, N5323, N5322, N5321,
		N5320, N5319}), .CI(1'b0), .SUM({ N5382, N5381, N5380, N5379, N5378,
		N5377, N5376, N5375, N5374, N5373, N5372, N5371, N5370, N5369, N5368,
		N5367, N5366, N5365, N5364, N5363, N5362, N5361, N5360, N5359, N5358,
		N5357, N5356, N5355, N5354, N5353, N5352, N5351}), .CO() );
	ID_DW01_add_32_2_test_1 sub_609 ( .A({ n331, n331, n331, n331, n331, n331,
		n331, n719, n695, n3990, n335, n336, n337, n878, n833, n340, IR_latched_15,
		IR_latched_14, IR_latched_13, IR_latched_12, IR_latched_11, IR_latched_10,
		IR_latched_9, IR_latched_8, n817, n3999, n888, IR_latched_4, IR_latched_3,
		IR_latched_2, IR_latched_1, IR_latched_0}), .B({ N5418, N5417, N5416,
		N5415, N5414, N5413, N5412, N5411, N5410, N5409, N5408, N5407, N5406,
		N5405, N5404, N5403, N5402, N5401, N5400, N5399, N5398, N5397, N5396,
		N5395, N5394, N5393, N5392, N5391, N5390, N5389, N5388, N5387}), .CI(1'b0),
		.SUM({ N5450, N5449, N5448, N5447, N5446, N5445, N5444, N5443, N5442,
		N5441, N5440, N5439, N5438, N5437, N5436, N5435, N5434, N5433, N5432,
		N5431, N5430, N5429, N5428, N5427, N5426, N5425, N5424, N5423, N5422,
		N5421, N5420, N5419}), .CO() );
	ID_DW01_add_32_1_test_1 sub_779 ( .A({ n887, n887, n887, n887, n887, n887,
		n887, n887, n887, n887, n887, n887, n887, n887, n887, n887, n887, IR_latched_14,
		IR_latched_13, IR_latched_12, IR_latched_11, IR_latched_10, n809, IR_latched_8,
		n817, n3999, n888, n831, IR_latched_3, IR_latched_2, IR_latched_1, IR_latched_0}),
		.B({ N6017, N6016, N6015, N6014, N6013, N6012, N6011, N6010, N6009, N6008,
		N6007, N6006, N6005, N6004, N6003, N6002, N6001, N6000, N5999, N5998,
		N5997, N5996, N5995, N5994, N5993, N5992, N5991, N5990, N5989, N5988,
		N5987, N5986}), .CI(1'b0), .SUM({ N6049, N6048, N6047, N6046, N6045,
		N6044, N6043, N6042, N6041, N6040, N6039, N6038, N6037, N6036, N6035,
		N6034, N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025,
		N6024, N6023, N6022, N6021, N6020, N6019, N6018}), .CO() );

endmodule


module IF_DW01_add_32_0_test_1 (  A, B, CI, SUM, CO );

input  CI;
input [31:0] A, B;
output  CO;
output [31:0] SUM;

wire A_0, A_1, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
	n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
	n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n49,
	n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
	n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
	n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
	n92, n93, n94, n95, n96, n97, n98, n99;

	assign A_1 = A[1];
	assign A_0 = A[0];
	assign SUM[1] = A_1;
	assign SUM[0] = A_0;

	nand2i_2 U10 ( .x(n72), .a(n106), .b(n107) );
	nand2i_4 U100 ( .x(n80), .a(n114), .b(n115) );
	exnor2_5 U101 ( .x(SUM[31]), .a(n82), .b(n121) );
	exnor2_5 U102 ( .x(SUM[30]), .a(n79), .b(n116) );
	exnor2_3 U103 ( .x(SUM[29]), .a(n122), .b(n81) );
	nand4_1 U104 ( .x(n94), .a(A[7]), .b(A[8]), .c(A[10]), .d(A[9]) );
	nand2_2 U106 ( .x(n111), .a(A[26]), .b(A[25]) );
	nand2_2 U107 ( .x(n114), .a(A[27]), .b(A[28]) );
	nand2_2 U108 ( .x(n83), .a(A[30]), .b(A[29]) );
	inv_5 U109 ( .x(n131), .a(n62) );
	nor2i_1 U11 ( .x(n71), .a(A[23]), .b(n72) );
	inv_5 U110 ( .x(n130), .a(n67) );
	inv_5 U111 ( .x(n129), .a(n72) );
	inv_5 U112 ( .x(n102), .a(n64) );
	inv_5 U113 ( .x(n107), .a(n69) );
	inv_5 U114 ( .x(n112), .a(n74) );
	inv_5 U115 ( .x(n115), .a(n77) );
	inv_6 U116 ( .x(n132), .a(n59) );
	nand2i_6 U117 ( .x(n64), .a(n99), .b(n131) );
	nand2i_6 U118 ( .x(n69), .a(n104), .b(n130) );
	nand2i_0 U119 ( .x(n109), .a(n128), .b(A[24]) );
	nor2_1 U12 ( .x(n68), .a(n69), .b(n70) );
	nand2_0 U120 ( .x(n106), .a(A[21]), .b(A[22]) );
	inv_0 U121 ( .x(n105), .a(A[22]) );
	nand2i_2 U13 ( .x(n59), .a(n94), .b(n92) );
	inv_2 U14 ( .x(n58), .a(n125) );
	nor2i_1 U15 ( .x(n57), .a(n58), .b(n59) );
	nand2i_2 U16 ( .x(n123), .a(n96), .b(n124) );
	nor2i_1 U17 ( .x(n49), .a(A[3]), .b(SUM[2]) );
	nand2i_2 U18 ( .x(n67), .a(n101), .b(n102) );
	nor2i_1 U19 ( .x(n66), .a(A[19]), .b(n67) );
	nor2_1 U20 ( .x(n63), .a(n64), .b(n65) );
	nand2i_2 U21 ( .x(n62), .a(n97), .b(n132) );
	inv_2 U22 ( .x(n61), .a(n126) );
	nor2i_1 U23 ( .x(n60), .a(n61), .b(n62) );
	inv_0 U24 ( .x(n125), .a(A[11]) );
	nand2i_2 U25 ( .x(n117), .a(n118), .b(n132) );
	inv_2 U26 ( .x(n92), .a(n53) );
	nand3i_1 U27 ( .x(n53), .a(SUM[2]), .b(n87), .c(n88) );
	nor2_1 U28 ( .x(n52), .a(n53), .b(n54) );
	nand2i_2 U29 ( .x(n56), .a(n91), .b(n92) );
	nand2i_2 U30 ( .x(n74), .a(n109), .b(n129) );
	nor2_1 U31 ( .x(n73), .a(n74), .b(n75) );
	nand2i_2 U32 ( .x(n77), .a(n111), .b(n112) );
	nor2_1 U33 ( .x(n76), .a(n77), .b(n78) );
	exnor2_1 U34 ( .x(SUM[24]), .a(n71), .b(n108) );
	exnor2_1 U35 ( .x(SUM[22]), .a(n68), .b(n105) );
	exnor2_1 U36 ( .x(SUM[12]), .a(n57), .b(n95) );
	exnor2_2 U37 ( .x(SUM[21]), .a(n107), .b(n70) );
	exnor2_2 U38 ( .x(SUM[25]), .a(n112), .b(n75) );
	exnor2_1 U39 ( .x(SUM[6]), .a(n50), .b(n86) );
	exnor2_1 U40 ( .x(SUM[4]), .a(n49), .b(n84) );
	inv_2 U41 ( .x(n120), .a(n51) );
	exnor2_1 U42 ( .x(SUM[11]), .a(n132), .b(n125) );
	exnor2_1 U43 ( .x(SUM[20]), .a(n66), .b(n103) );
	exnor2_3 U44 ( .x(SUM[23]), .a(n129), .b(n128) );
	exnor2_1 U45 ( .x(SUM[18]), .a(n63), .b(n100) );
	exnor2_1 U46 ( .x(SUM[17]), .a(n102), .b(n65) );
	exnor2_1 U47 ( .x(SUM[15]), .a(n131), .b(n126) );
	exnor2_1 U48 ( .x(SUM[16]), .a(n60), .b(n98) );
	exnor2_1 U49 ( .x(SUM[13]), .a(n124), .b(n96) );
	nand2i_2 U5 ( .x(n104), .a(n127), .b(A[20]) );
	inv_2 U50 ( .x(n124), .a(n117) );
	exnor2_2 U51 ( .x(SUM[19]), .a(n130), .b(n127) );
	exnor2_2 U52 ( .x(SUM[7]), .a(n92), .b(n54) );
	inv_2 U53 ( .x(n54), .a(A[7]) );
	exnor2_1 U54 ( .x(SUM[9]), .a(n119), .b(n90) );
	inv_2 U55 ( .x(n119), .a(n56) );
	exnor2_1 U56 ( .x(SUM[8]), .a(n52), .b(n89) );
	exnor2_1 U57 ( .x(SUM[10]), .a(n55), .b(n93) );
	exor2_1 U58 ( .x(SUM[3]), .a(A[3]), .b(A[2]) );
	inv_2 U59 ( .x(SUM[2]), .a(A[2]) );
	nand2i_0 U6 ( .x(n99), .a(n126), .b(A[16]) );
	inv_1 U60 ( .x(n103), .a(A[20]) );
	inv_0 U61 ( .x(n75), .a(A[25]) );
	inv_2 U62 ( .x(n81), .a(A[29]) );
	exnor2_1 U63 ( .x(SUM[26]), .a(n73), .b(n110) );
	exnor2_1 U64 ( .x(SUM[27]), .a(n115), .b(n78) );
	exnor2_1 U65 ( .x(SUM[28]), .a(n76), .b(n113) );
	inv_2 U66 ( .x(n122), .a(n80) );
	inv_0 U67 ( .x(n108), .a(A[24]) );
	inv_0 U69 ( .x(n70), .a(A[21]) );
	nor2i_1 U7 ( .x(n88), .a(A[3]), .b(n84) );
	inv_0 U70 ( .x(n127), .a(A[19]) );
	inv_2 U71 ( .x(n78), .a(A[27]) );
	inv_2 U72 ( .x(n113), .a(A[28]) );
	inv_2 U73 ( .x(n116), .a(A[30]) );
	inv_2 U74 ( .x(n121), .a(A[31]) );
	inv_2 U75 ( .x(n128), .a(A[23]) );
	exnor2_1 U76 ( .x(SUM[5]), .a(n120), .b(n85) );
	inv_0 U77 ( .x(n98), .a(A[16]) );
	inv_0 U78 ( .x(n126), .a(A[15]) );
	inv_0 U79 ( .x(n65), .a(A[17]) );
	inv_0 U80 ( .x(n89), .a(A[8]) );
	nor2i_0 U81 ( .x(n87), .a(A[6]), .b(n85) );
	inv_0 U82 ( .x(n86), .a(A[6]) );
	inv_0 U83 ( .x(n96), .a(A[13]) );
	nand2_0 U84 ( .x(n101), .a(A[17]), .b(A[18]) );
	inv_0 U85 ( .x(n100), .a(A[18]) );
	nand3i_0 U86 ( .x(n51), .a(SUM[2]), .b(A[4]), .c(A[3]) );
	inv_1 U87 ( .x(n84), .a(A[4]) );
	exnor2_1 U88 ( .x(SUM[14]), .a(A[14]), .b(n123) );
	inv_0 U89 ( .x(n93), .a(A[10]) );
	inv_0 U9 ( .x(n110), .a(A[26]) );
	inv_0 U90 ( .x(n90), .a(A[9]) );
	nor2i_0 U91 ( .x(n55), .a(A[9]), .b(n56) );
	nand2_0 U92 ( .x(n91), .a(A[7]), .b(A[8]) );
	inv_0 U93 ( .x(n95), .a(A[12]) );
	nand2i_0 U94 ( .x(n118), .a(n125), .b(A[12]) );
	nand4i_1 U95 ( .x(n97), .a(n125), .b(A[13]), .c(A[12]), .d(A[14]) );
	nor2i_0 U96 ( .x(n50), .a(A[5]), .b(n51) );
	inv_0 U97 ( .x(n85), .a(A[5]) );
	nor2_5 U98 ( .x(n79), .a(n80), .b(n81) );
	nor2_5 U99 ( .x(n82), .a(n80), .b(n83) );

endmodule


module IF_test_1_desync (  NPC, PC, IR_latched, reset, branch_sig, branch_address,
	IR, stall, counter, test_si1, test_so1, test_si2, test_se, sync_sel, global_g1,
	global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );

input  reset, branch_sig, stall, test_si1, test_si2, test_se, sync_sel,
	global_g1, global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
input [1:0] counter;
input [31:0] branch_address, IR;
output  test_so1;
output [31:0] NPC, PC, IR_latched;

wire IR_curr_0, IR_curr_1, IR_curr_10, IR_curr_11, IR_curr_12, IR_curr_13,
	IR_curr_14, IR_curr_15, IR_curr_16, IR_curr_17, IR_curr_18, IR_curr_19,
	IR_curr_2, IR_curr_20, IR_curr_21, IR_curr_22, IR_curr_23, IR_curr_24,
	IR_curr_25, IR_curr_26, IR_curr_27, IR_curr_28, IR_curr_29, IR_curr_3,
	IR_curr_30, IR_curr_31, IR_curr_4, IR_curr_5, IR_curr_6, IR_curr_7, IR_curr_8,
	IR_curr_9, IR_curr_reg_0__m2s, IR_curr_reg_10__m2s, IR_curr_reg_11__m2s,
	IR_curr_reg_12__m2s, IR_curr_reg_13__m2s, IR_curr_reg_14__m2s, IR_curr_reg_15__m2s,
	IR_curr_reg_16__m2s, IR_curr_reg_17__m2s, IR_curr_reg_18__m2s, IR_curr_reg_19__m2s,
	IR_curr_reg_1__m2s, IR_curr_reg_20__m2s, IR_curr_reg_21__m2s, IR_curr_reg_22__m2s,
	IR_curr_reg_23__m2s, IR_curr_reg_24__m2s, IR_curr_reg_25__m2s, IR_curr_reg_26__m2s,
	IR_curr_reg_27__m2s, IR_curr_reg_28__m2s, IR_curr_reg_29__m2s, IR_curr_reg_2__m2s,
	IR_curr_reg_30__m2s, IR_curr_reg_31__m2s, IR_curr_reg_3__m2s, IR_curr_reg_4__m2s,
	IR_curr_reg_5__m2s, IR_curr_reg_6__m2s, IR_curr_reg_7__m2s, IR_curr_reg_8__m2s,
	IR_curr_reg_9__m2s, IR_latched_reg_0__m2s, IR_latched_reg_10__m2s, IR_latched_reg_11__m2s,
	IR_latched_reg_12__m2s, IR_latched_reg_13__m2s, IR_latched_reg_14__m2s,
	IR_latched_reg_15__m2s, IR_latched_reg_16__m2s, IR_latched_reg_17__m2s,
	IR_latched_reg_18__m2s, IR_latched_reg_19__m2s, IR_latched_reg_1__m2s,
	IR_latched_reg_20__m2s, IR_latched_reg_21__m2s, IR_latched_reg_22__m2s,
	IR_latched_reg_23__m2s, IR_latched_reg_24__m2s, IR_latched_reg_25__m2s,
	IR_latched_reg_26__m2s, IR_latched_reg_27__m2s, IR_latched_reg_28__m2s,
	IR_latched_reg_29__m2s, IR_latched_reg_2__m2s, IR_latched_reg_30__m2s,
	IR_latched_reg_31__m2s, IR_latched_reg_3__m2s, IR_latched_reg_4__m2s,
	IR_latched_reg_5__m2s, IR_latched_reg_6__m2s, IR_latched_reg_7__m2s, IR_latched_reg_8__m2s,
	IR_latched_reg_9__m2s, IR_previous_0, IR_previous_1, IR_previous_10, IR_previous_11,
	IR_previous_12, IR_previous_13, IR_previous_14, IR_previous_15, IR_previous_16,
	IR_previous_17, IR_previous_18, IR_previous_19, IR_previous_2, IR_previous_20,
	IR_previous_21, IR_previous_22, IR_previous_23, IR_previous_24, IR_previous_25,
	IR_previous_26, IR_previous_27, IR_previous_28, IR_previous_29, IR_previous_3,
	IR_previous_30, IR_previous_31, IR_previous_4, IR_previous_5, IR_previous_6,
	IR_previous_7, IR_previous_8, IR_previous_9, IR_previous_reg_0__m2s, IR_previous_reg_10__m2s,
	IR_previous_reg_11__m2s, IR_previous_reg_12__m2s, IR_previous_reg_13__m2s,
	IR_previous_reg_14__m2s, IR_previous_reg_15__m2s, IR_previous_reg_16__m2s,
	IR_previous_reg_17__m2s, IR_previous_reg_18__m2s, IR_previous_reg_19__m2s,
	IR_previous_reg_1__m2s, IR_previous_reg_20__m2s, IR_previous_reg_21__m2s,
	IR_previous_reg_22__m2s, IR_previous_reg_23__m2s, IR_previous_reg_24__m2s,
	IR_previous_reg_25__m2s, IR_previous_reg_26__m2s, IR_previous_reg_27__m2s,
	IR_previous_reg_28__m2s, IR_previous_reg_29__m2s, IR_previous_reg_2__m2s,
	IR_previous_reg_30__m2s, IR_previous_reg_31__m2s, IR_previous_reg_3__m2s,
	IR_previous_reg_4__m2s, IR_previous_reg_5__m2s, IR_previous_reg_6__m2s,
	IR_previous_reg_7__m2s, IR_previous_reg_8__m2s, IR_previous_reg_9__m2s,
	N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
	N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
	N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135,
	N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147,
	N148, N149, N150, N152, N17, N18, N19, N20, N21, N215, N22, N23, N24,
	N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38,
	N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N50, N87, N88, N89,
	N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, NPC_reg_0__m2s, NPC_reg_10__m2s,
	NPC_reg_11__m2s, NPC_reg_12__m2s, NPC_reg_13__m2s, NPC_reg_14__m2s, NPC_reg_15__m2s,
	NPC_reg_16__m2s, NPC_reg_17__m2s, NPC_reg_18__m2s, NPC_reg_19__m2s, NPC_reg_1__m2s,
	NPC_reg_20__m2s, NPC_reg_21__m2s, NPC_reg_22__m2s, NPC_reg_23__m2s, NPC_reg_24__m2s,
	NPC_reg_25__m2s, NPC_reg_26__m2s, NPC_reg_27__m2s, NPC_reg_28__m2s, NPC_reg_29__m2s,
	NPC_reg_2__m2s, NPC_reg_30__m2s, NPC_reg_31__m2s, NPC_reg_3__m2s, NPC_reg_4__m2s,
	NPC_reg_5__m2s, NPC_reg_6__m2s, NPC_reg_7__m2s, NPC_reg_8__m2s, NPC_reg_9__m2s,
	PC_reg_0__m2s, PC_reg_10__m2s, PC_reg_11__m2s, PC_reg_12__m2s, PC_reg_13__m2s,
	PC_reg_14__m2s, PC_reg_15__m2s, PC_reg_16__m2s, PC_reg_17__m2s, PC_reg_18__m2s,
	PC_reg_19__m2s, PC_reg_1__m2s, PC_reg_20__m2s, PC_reg_21__m2s, PC_reg_22__m2s,
	PC_reg_23__m2s, PC_reg_24__m2s, PC_reg_25__m2s, PC_reg_26__m2s, PC_reg_27__m2s,
	PC_reg_28__m2s, PC_reg_29__m2s, PC_reg_2__m2s, PC_reg_30__m2s, PC_reg_31__m2s,
	PC_reg_3__m2s, PC_reg_4__m2s, PC_reg_5__m2s, PC_reg_6__m2s, PC_reg_7__m2s,
	PC_reg_8__m2s, PC_reg_9__m2s, n10, n100, n101, n102, n104, n105, n106,
	n107, n108, n109, n11, n110, n111, n112, n113, n114, n115, n116, n117,
	n118, n119, n12, n120, n121, n122, n123, n124, n125, n126, n127, n128,
	n129, n13, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
	n14, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n15,
	n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n16, n160,
	n161, n162, n163, n164, n165, n166, n167, n168, n169, n17, n170, n171,
	n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
	n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
	n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
	n208, n209, n210, n211, n212, n213, n214, n215, n217, n218, n22, n221,
	n222, n223, n224, n225, n226, n227, n228, n229, n23, n230, n231, n232,
	n233, n234, n235, n236, n237, n238, n239, n24, n240, n241, n242, n243,
	n244, n245, n246, n247, n248, n249, n25, n250, n251, n252, n253, n254,
	n255, n256, n257, n258, n259, n26, n260, n261, n262, n263, n264, n265,
	n266, n267, n268, n269, n27, n270, n271, n272, n273, n274, n275, n276,
	n277, n278, n279, n28, n280, n281, n282, n283, n284, n285, n286, n287,
	n288, n289, n29, n290, n291, n292, n293, n294, n295, n296, n297, n298,
	n299, n30, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
	n31, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n32,
	n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n33, n330,
	n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
	n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
	n355, n356, n357, n358, n36, n360, n37, n38, n39, n4, n40, n41, n42, n43,
	n44, n45, n46, n47, n48, n49, n5, n50, n51, n52, n53, n54, n55, n56, n57,
	n58, n59, n6, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n7, n70,
	n71, n72, n73, n74, n75, n76, n77, n78, n79, n8, n80, n81, n82, n83, n84,
	n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
	n99, stalled_reg__m2s;


	smlatnr_1 IR_curr_reg_0__master ( .q(IR_curr_reg_0__m2s), .qb(), .d(n136),
		.sdi(test_si1), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_0__slave ( .q(IR_curr_0), .qb(n358), .d(IR_curr_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_10__master ( .q(IR_curr_reg_10__m2s), .qb(), .d(n146),
		.sdi(n349), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_10__slave ( .q(IR_curr_10), .qb(n348), .d(IR_curr_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_11__master ( .q(IR_curr_reg_11__m2s), .qb(), .d(n147),
		.sdi(n348), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_11__slave ( .q(IR_curr_11), .qb(n347), .d(IR_curr_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_12__master ( .q(IR_curr_reg_12__m2s), .qb(), .d(n148),
		.sdi(n347), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_12__slave ( .q(IR_curr_12), .qb(n346), .d(IR_curr_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_13__master ( .q(IR_curr_reg_13__m2s), .qb(), .d(n149),
		.sdi(n346), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_13__slave ( .q(IR_curr_13), .qb(n345), .d(IR_curr_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_14__master ( .q(IR_curr_reg_14__m2s), .qb(), .d(n150),
		.sdi(n345), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_14__slave ( .q(IR_curr_14), .qb(n344), .d(IR_curr_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_15__master ( .q(IR_curr_reg_15__m2s), .qb(), .d(n151),
		.sdi(n344), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_15__slave ( .q(IR_curr_15), .qb(n343), .d(IR_curr_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_16__master ( .q(IR_curr_reg_16__m2s), .qb(), .d(n152),
		.sdi(n343), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_16__slave ( .q(IR_curr_16), .qb(n342), .d(IR_curr_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_17__master ( .q(IR_curr_reg_17__m2s), .qb(), .d(n153),
		.sdi(n342), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_17__slave ( .q(IR_curr_17), .qb(n341), .d(IR_curr_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_18__master ( .q(IR_curr_reg_18__m2s), .qb(), .d(n154),
		.sdi(n341), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_18__slave ( .q(IR_curr_18), .qb(n340), .d(IR_curr_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_19__master ( .q(IR_curr_reg_19__m2s), .qb(), .d(n155),
		.sdi(n340), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_19__slave ( .q(IR_curr_19), .qb(n339), .d(IR_curr_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_1__master ( .q(IR_curr_reg_1__m2s), .qb(), .d(n137),
		.sdi(n358), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_1__slave ( .q(IR_curr_1), .qb(n357), .d(IR_curr_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_20__master ( .q(IR_curr_reg_20__m2s), .qb(), .d(n156),
		.sdi(n339), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_20__slave ( .q(IR_curr_20), .qb(n338), .d(IR_curr_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_21__master ( .q(IR_curr_reg_21__m2s), .qb(), .d(n157),
		.sdi(n338), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_21__slave ( .q(IR_curr_21), .qb(n337), .d(IR_curr_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_22__master ( .q(IR_curr_reg_22__m2s), .qb(), .d(n158),
		.sdi(n337), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_22__slave ( .q(IR_curr_22), .qb(n336), .d(IR_curr_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_23__master ( .q(IR_curr_reg_23__m2s), .qb(), .d(n159),
		.sdi(n336), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_23__slave ( .q(IR_curr_23), .qb(n335), .d(IR_curr_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_24__master ( .q(IR_curr_reg_24__m2s), .qb(), .d(n160),
		.sdi(n335), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_24__slave ( .q(IR_curr_24), .qb(n334), .d(IR_curr_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_25__master ( .q(IR_curr_reg_25__m2s), .qb(), .d(n161),
		.sdi(n334), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_25__slave ( .q(IR_curr_25), .qb(n333), .d(IR_curr_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_26__master ( .q(IR_curr_reg_26__m2s), .qb(), .d(n162),
		.sdi(n333), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_26__slave ( .q(IR_curr_26), .qb(n332), .d(IR_curr_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_27__master ( .q(IR_curr_reg_27__m2s), .qb(), .d(n163),
		.sdi(n332), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_27__slave ( .q(IR_curr_27), .qb(n331), .d(IR_curr_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_28__master ( .q(IR_curr_reg_28__m2s), .qb(), .d(n164),
		.sdi(n331), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_28__slave ( .q(IR_curr_28), .qb(n330), .d(IR_curr_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_29__master ( .q(IR_curr_reg_29__m2s), .qb(), .d(n165),
		.sdi(n330), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_29__slave ( .q(IR_curr_29), .qb(n329), .d(IR_curr_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_2__master ( .q(IR_curr_reg_2__m2s), .qb(), .d(n138),
		.sdi(n357), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_2__slave ( .q(IR_curr_2), .qb(n356), .d(IR_curr_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_30__master ( .q(IR_curr_reg_30__m2s), .qb(), .d(n166),
		.sdi(n329), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_30__slave ( .q(IR_curr_30), .qb(n328), .d(IR_curr_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_31__master ( .q(IR_curr_reg_31__m2s), .qb(), .d(n167),
		.sdi(n328), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_31__slave ( .q(IR_curr_31), .qb(n327), .d(IR_curr_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_3__master ( .q(IR_curr_reg_3__m2s), .qb(), .d(n139),
		.sdi(n356), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_3__slave ( .q(IR_curr_3), .qb(n355), .d(IR_curr_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_4__master ( .q(IR_curr_reg_4__m2s), .qb(), .d(n140),
		.sdi(n355), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_4__slave ( .q(IR_curr_4), .qb(n354), .d(IR_curr_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_5__master ( .q(IR_curr_reg_5__m2s), .qb(), .d(n141),
		.sdi(n354), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n41), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_5__slave ( .q(IR_curr_5), .qb(n353), .d(IR_curr_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n41), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_6__master ( .q(IR_curr_reg_6__m2s), .qb(), .d(n142),
		.sdi(n353), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_6__slave ( .q(IR_curr_6), .qb(n352), .d(IR_curr_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_7__master ( .q(IR_curr_reg_7__m2s), .qb(), .d(n143),
		.sdi(n352), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_7__slave ( .q(IR_curr_7), .qb(n351), .d(IR_curr_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_8__master ( .q(IR_curr_reg_8__m2s), .qb(), .d(n144),
		.sdi(n351), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_8__slave ( .q(IR_curr_8), .qb(n350), .d(IR_curr_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_curr_reg_9__master ( .q(IR_curr_reg_9__m2s), .qb(), .d(n145),
		.sdi(n350), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 IR_curr_reg_9__slave ( .q(IR_curr_9), .qb(n349), .d(IR_curr_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_0__master ( .q(IR_latched_reg_0__m2s), .qb(),
		.d(N119), .sdi(n327), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_0__slave ( .q(IR_latched[0]), .qb(n326), .d(IR_latched_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_10__master ( .q(IR_latched_reg_10__m2s), .qb(),
		.d(N129), .sdi(n317), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_10__slave ( .q(IR_latched[10]), .qb(n316), .d(IR_latched_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_11__master ( .q(IR_latched_reg_11__m2s), .qb(),
		.d(N130), .sdi(n316), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_11__slave ( .q(IR_latched[11]), .qb(n315), .d(IR_latched_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_12__master ( .q(IR_latched_reg_12__m2s), .qb(),
		.d(N131), .sdi(n315), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_12__slave ( .q(IR_latched[12]), .qb(n314), .d(IR_latched_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_13__master ( .q(IR_latched_reg_13__m2s), .qb(),
		.d(N132), .sdi(n314), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_13__slave ( .q(IR_latched[13]), .qb(n313), .d(IR_latched_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_14__master ( .q(IR_latched_reg_14__m2s), .qb(),
		.d(N133), .sdi(n313), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_14__slave ( .q(IR_latched[14]), .qb(n312), .d(IR_latched_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_15__master ( .q(IR_latched_reg_15__m2s), .qb(),
		.d(N134), .sdi(n312), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_15__slave ( .q(IR_latched[15]), .qb(n311), .d(IR_latched_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_16__master ( .q(IR_latched_reg_16__m2s), .qb(),
		.d(N135), .sdi(n311), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_16__slave ( .q(IR_latched[16]), .qb(n310), .d(IR_latched_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_17__master ( .q(IR_latched_reg_17__m2s), .qb(),
		.d(N136), .sdi(n310), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_17__slave ( .q(IR_latched[17]), .qb(n309), .d(IR_latched_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_18__master ( .q(IR_latched_reg_18__m2s), .qb(),
		.d(N137), .sdi(n309), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_18__slave ( .q(IR_latched[18]), .qb(n308), .d(IR_latched_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_19__master ( .q(IR_latched_reg_19__m2s), .qb(),
		.d(N138), .sdi(n308), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_19__slave ( .q(IR_latched[19]), .qb(n307), .d(IR_latched_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_1__master ( .q(IR_latched_reg_1__m2s), .qb(),
		.d(N120), .sdi(n326), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_1__slave ( .q(IR_latched[1]), .qb(n325), .d(IR_latched_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_20__master ( .q(IR_latched_reg_20__m2s), .qb(),
		.d(N139), .sdi(n307), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_20__slave ( .q(IR_latched[20]), .qb(n306), .d(IR_latched_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_21__master ( .q(IR_latched_reg_21__m2s), .qb(),
		.d(N140), .sdi(n306), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_21__slave ( .q(IR_latched[21]), .qb(n305), .d(IR_latched_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_22__master ( .q(IR_latched_reg_22__m2s), .qb(),
		.d(N141), .sdi(n305), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_22__slave ( .q(IR_latched[22]), .qb(n304), .d(IR_latched_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_23__master ( .q(IR_latched_reg_23__m2s), .qb(),
		.d(N142), .sdi(n304), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_23__slave ( .q(IR_latched[23]), .qb(n303), .d(IR_latched_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_24__master ( .q(IR_latched_reg_24__m2s), .qb(),
		.d(N143), .sdi(n303), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_24__slave ( .q(IR_latched[24]), .qb(n302), .d(IR_latched_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_25__master ( .q(IR_latched_reg_25__m2s), .qb(),
		.d(N144), .sdi(n302), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_25__slave ( .q(IR_latched[25]), .qb(n301), .d(IR_latched_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_26__master ( .q(IR_latched_reg_26__m2s), .qb(),
		.d(N145), .sdi(n301), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_26__slave ( .q(IR_latched[26]), .qb(n300), .d(IR_latched_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_27__master ( .q(IR_latched_reg_27__m2s), .qb(),
		.d(N146), .sdi(n300), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_27__slave ( .q(IR_latched[27]), .qb(n299), .d(IR_latched_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_28__master ( .q(IR_latched_reg_28__m2s), .qb(),
		.d(N147), .sdi(n299), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_28__slave ( .q(IR_latched[28]), .qb(n298), .d(IR_latched_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_29__master ( .q(IR_latched_reg_29__m2s), .qb(),
		.d(N148), .sdi(n298), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_29__slave ( .q(IR_latched[29]), .qb(n297), .d(IR_latched_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_2__master ( .q(IR_latched_reg_2__m2s), .qb(),
		.d(N121), .sdi(n325), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_2__slave ( .q(IR_latched[2]), .qb(n324), .d(IR_latched_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_30__master ( .q(IR_latched_reg_30__m2s), .qb(),
		.d(N149), .sdi(n297), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_30__slave ( .q(IR_latched[30]), .qb(n296), .d(IR_latched_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_31__master ( .q(IR_latched_reg_31__m2s), .qb(),
		.d(N150), .sdi(n296), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n37),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_31__slave ( .q(IR_latched[31]), .qb(n295), .d(IR_latched_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n37), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_3__master ( .q(IR_latched_reg_3__m2s), .qb(),
		.d(N122), .sdi(n324), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_3__slave ( .q(IR_latched[3]), .qb(n323), .d(IR_latched_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_4__master ( .q(IR_latched_reg_4__m2s), .qb(),
		.d(N123), .sdi(n323), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_4__slave ( .q(IR_latched[4]), .qb(n322), .d(IR_latched_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_5__master ( .q(IR_latched_reg_5__m2s), .qb(),
		.d(N124), .sdi(n322), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_5__slave ( .q(IR_latched[5]), .qb(n321), .d(IR_latched_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_6__master ( .q(IR_latched_reg_6__m2s), .qb(),
		.d(N125), .sdi(n321), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_6__slave ( .q(IR_latched[6]), .qb(n320), .d(IR_latched_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_7__master ( .q(IR_latched_reg_7__m2s), .qb(),
		.d(N126), .sdi(n320), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_7__slave ( .q(IR_latched[7]), .qb(n319), .d(IR_latched_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_8__master ( .q(IR_latched_reg_8__m2s), .qb(),
		.d(N127), .sdi(n319), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_8__slave ( .q(IR_latched[8]), .qb(n318), .d(IR_latched_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_latched_reg_9__master ( .q(IR_latched_reg_9__m2s), .qb(),
		.d(N128), .sdi(n318), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_latched_reg_9__slave ( .q(IR_latched[9]), .qb(n317), .d(IR_latched_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_0__master ( .q(IR_previous_reg_0__m2s), .qb(),
		.d(n104), .sdi(n295), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_0__slave ( .q(IR_previous_0), .qb(n294), .d(IR_previous_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_10__master ( .q(IR_previous_reg_10__m2s), .qb(),
		.d(n114), .sdi(n285), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_10__slave ( .q(IR_previous_10), .qb(n284), .d(IR_previous_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_11__master ( .q(IR_previous_reg_11__m2s), .qb(),
		.d(n115), .sdi(n284), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_11__slave ( .q(IR_previous_11), .qb(n283), .d(IR_previous_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_12__master ( .q(IR_previous_reg_12__m2s), .qb(),
		.d(n116), .sdi(n283), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_12__slave ( .q(IR_previous_12), .qb(n282), .d(IR_previous_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_13__master ( .q(IR_previous_reg_13__m2s), .qb(),
		.d(n117), .sdi(n282), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_13__slave ( .q(IR_previous_13), .qb(n281), .d(IR_previous_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_14__master ( .q(IR_previous_reg_14__m2s), .qb(),
		.d(n118), .sdi(n281), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n42),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_14__slave ( .q(IR_previous_14), .qb(n280), .d(IR_previous_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n42), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_15__master ( .q(IR_previous_reg_15__m2s), .qb(),
		.d(n119), .sdi(n280), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_15__slave ( .q(IR_previous_15), .qb(n279), .d(IR_previous_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_16__master ( .q(IR_previous_reg_16__m2s), .qb(),
		.d(n120), .sdi(n279), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_16__slave ( .q(IR_previous_16), .qb(n278), .d(IR_previous_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_17__master ( .q(IR_previous_reg_17__m2s), .qb(),
		.d(n121), .sdi(n278), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_17__slave ( .q(IR_previous_17), .qb(n277), .d(IR_previous_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_18__master ( .q(IR_previous_reg_18__m2s), .qb(),
		.d(n122), .sdi(n277), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_18__slave ( .q(IR_previous_18), .qb(n276), .d(IR_previous_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_19__master ( .q(IR_previous_reg_19__m2s), .qb(),
		.d(n123), .sdi(n276), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_19__slave ( .q(IR_previous_19), .qb(n275), .d(IR_previous_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_1__master ( .q(IR_previous_reg_1__m2s), .qb(),
		.d(n105), .sdi(n294), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_1__slave ( .q(IR_previous_1), .qb(n293), .d(IR_previous_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_20__master ( .q(IR_previous_reg_20__m2s), .qb(),
		.d(n124), .sdi(n275), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_20__slave ( .q(IR_previous_20), .qb(n274), .d(IR_previous_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_21__master ( .q(IR_previous_reg_21__m2s), .qb(),
		.d(n125), .sdi(n274), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_21__slave ( .q(IR_previous_21), .qb(n273), .d(IR_previous_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_22__master ( .q(IR_previous_reg_22__m2s), .qb(),
		.d(n126), .sdi(n273), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_22__slave ( .q(IR_previous_22), .qb(n272), .d(IR_previous_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_23__master ( .q(IR_previous_reg_23__m2s), .qb(),
		.d(n127), .sdi(n272), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_23__slave ( .q(IR_previous_23), .qb(n271), .d(IR_previous_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_24__master ( .q(IR_previous_reg_24__m2s), .qb(),
		.d(n128), .sdi(n271), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_24__slave ( .q(IR_previous_24), .qb(n270), .d(IR_previous_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_25__master ( .q(IR_previous_reg_25__m2s), .qb(),
		.d(n129), .sdi(n270), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_25__slave ( .q(IR_previous_25), .qb(n269), .d(IR_previous_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_26__master ( .q(IR_previous_reg_26__m2s), .qb(),
		.d(n130), .sdi(n269), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_26__slave ( .q(IR_previous_26), .qb(n268), .d(IR_previous_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_27__master ( .q(IR_previous_reg_27__m2s), .qb(),
		.d(n131), .sdi(n268), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_27__slave ( .q(IR_previous_27), .qb(n267), .d(IR_previous_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_28__master ( .q(IR_previous_reg_28__m2s), .qb(),
		.d(n132), .sdi(n267), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_28__slave ( .q(IR_previous_28), .qb(n266), .d(IR_previous_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_29__master ( .q(IR_previous_reg_29__m2s), .qb(),
		.d(n133), .sdi(n266), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_29__slave ( .q(IR_previous_29), .qb(n265), .d(IR_previous_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_2__master ( .q(IR_previous_reg_2__m2s), .qb(),
		.d(n106), .sdi(n293), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_2__slave ( .q(IR_previous_2), .qb(n292), .d(IR_previous_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_30__master ( .q(IR_previous_reg_30__m2s), .qb(),
		.d(n134), .sdi(n265), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_30__slave ( .q(IR_previous_30), .qb(n264), .d(IR_previous_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_31__master ( .q(IR_previous_reg_31__m2s), .qb(),
		.d(n135), .sdi(n264), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_31__slave ( .q(IR_previous_31), .qb(n263), .d(IR_previous_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_3__master ( .q(IR_previous_reg_3__m2s), .qb(),
		.d(n107), .sdi(n292), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_3__slave ( .q(IR_previous_3), .qb(n291), .d(IR_previous_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_4__master ( .q(IR_previous_reg_4__m2s), .qb(),
		.d(n108), .sdi(n291), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_4__slave ( .q(IR_previous_4), .qb(n290), .d(IR_previous_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_5__master ( .q(IR_previous_reg_5__m2s), .qb(),
		.d(n109), .sdi(n290), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_5__slave ( .q(IR_previous_5), .qb(n289), .d(IR_previous_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_6__master ( .q(IR_previous_reg_6__m2s), .qb(),
		.d(n110), .sdi(n289), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_6__slave ( .q(IR_previous_6), .qb(n288), .d(IR_previous_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_7__master ( .q(IR_previous_reg_7__m2s), .qb(),
		.d(n111), .sdi(n288), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_7__slave ( .q(IR_previous_7), .qb(n287), .d(IR_previous_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_8__master ( .q(IR_previous_reg_8__m2s), .qb(),
		.d(n112), .sdi(n287), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_8__slave ( .q(IR_previous_8), .qb(n286), .d(IR_previous_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 IR_previous_reg_9__master ( .q(IR_previous_reg_9__m2s), .qb(),
		.d(n113), .sdi(n286), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 IR_previous_reg_9__slave ( .q(IR_previous_9), .qb(n285), .d(IR_previous_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_0__master ( .q(NPC_reg_0__m2s), .qb(), .d(N87), .sdi(n263),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_0__slave ( .q(NPC[0]), .qb(n262), .d(NPC_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_10__master ( .q(NPC_reg_10__m2s), .qb(), .d(N97), .sdi(n22),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_10__slave ( .q(NPC[10]), .qb(n24), .d(NPC_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_11__master ( .q(NPC_reg_11__m2s), .qb(), .d(N98), .sdi(n24),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_11__slave ( .q(n205), .qb(n257), .d(NPC_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_12__master ( .q(NPC_reg_12__m2s), .qb(), .d(N99), .sdi(n257),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_12__slave ( .q(NPC[12]), .qb(n28), .d(NPC_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_13__master ( .q(NPC_reg_13__m2s), .qb(), .d(N100), .sdi(n28),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_13__slave ( .q(NPC[13]), .qb(n14), .d(NPC_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_14__master ( .q(NPC_reg_14__m2s), .qb(), .d(N101), .sdi(n14),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_14__slave ( .q(n360), .qb(n12), .d(NPC_reg_14__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_15__master ( .q(NPC_reg_15__m2s), .qb(), .d(N102), .sdi(n12),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_15__slave ( .q(n204), .qb(n256), .d(NPC_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_16__master ( .q(NPC_reg_16__m2s), .qb(), .d(N103), .sdi(n256),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_16__slave ( .q(NPC[16]), .qb(n255), .d(NPC_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_17__master ( .q(NPC_reg_17__m2s), .qb(), .d(N104), .sdi(n255),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_17__slave ( .q(NPC[17]), .qb(n10), .d(NPC_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_18__master ( .q(NPC_reg_18__m2s), .qb(), .d(N105), .sdi(n10),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_18__slave ( .q(NPC[18]), .qb(n254), .d(NPC_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_19__master ( .q(NPC_reg_19__m2s), .qb(), .d(N106), .sdi(n254),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_19__slave ( .q(NPC[19]), .qb(n253), .d(NPC_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_1__master ( .q(NPC_reg_1__m2s), .qb(), .d(N88), .sdi(n262),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_1__slave ( .q(NPC[1]), .qb(n261), .d(NPC_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_20__master ( .q(NPC_reg_20__m2s), .qb(), .d(N107), .sdi(n253),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_20__slave ( .q(NPC[20]), .qb(n252), .d(NPC_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_21__master ( .q(NPC_reg_21__m2s), .qb(), .d(N108), .sdi(n252),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_21__slave ( .q(NPC[21]), .qb(n251), .d(NPC_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_22__master ( .q(NPC_reg_22__m2s), .qb(), .d(N109), .sdi(n251),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_22__slave ( .q(NPC[22]), .qb(n250), .d(NPC_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_23__master ( .q(NPC_reg_23__m2s), .qb(), .d(N110), .sdi(n250),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_23__slave ( .q(NPC[23]), .qb(n249), .d(NPC_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_24__master ( .q(NPC_reg_24__m2s), .qb(), .d(N111), .sdi(n249),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n91), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_24__slave ( .q(NPC[24]), .qb(n248), .d(NPC_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n91), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_25__master ( .q(NPC_reg_25__m2s), .qb(), .d(N112), .sdi(n248),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_25__slave ( .q(NPC[25]), .qb(n247), .d(NPC_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_26__master ( .q(NPC_reg_26__m2s), .qb(), .d(N113), .sdi(n247),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_26__slave ( .q(NPC[26]), .qb(n246), .d(NPC_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_27__master ( .q(NPC_reg_27__m2s), .qb(), .d(N114), .sdi(n246),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_27__slave ( .q(NPC[27]), .qb(n245), .d(NPC_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_28__master ( .q(NPC_reg_28__m2s), .qb(), .d(N115), .sdi(n245),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_28__slave ( .q(NPC[28]), .qb(n244), .d(NPC_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_29__master ( .q(NPC_reg_29__m2s), .qb(), .d(N116), .sdi(n244),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_29__slave ( .q(NPC[29]), .qb(n243), .d(NPC_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_2__master ( .q(NPC_reg_2__m2s), .qb(), .d(N89), .sdi(n261),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_2__slave ( .q(n210), .qb(n32), .d(NPC_reg_2__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_30__master ( .q(NPC_reg_30__m2s), .qb(), .d(N117), .sdi(n243),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_30__slave ( .q(NPC[30]), .qb(n242), .d(NPC_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_31__master ( .q(NPC_reg_31__m2s), .qb(), .d(N118), .sdi(test_si2),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_31__slave ( .q(NPC[31]), .qb(), .d(NPC_reg_31__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_3__master ( .q(NPC_reg_3__m2s), .qb(), .d(N90), .sdi(n32),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_3__slave ( .q(n209), .qb(n30), .d(NPC_reg_3__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_4__master ( .q(NPC_reg_4__m2s), .qb(), .d(N91), .sdi(n30),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n40), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 NPC_reg_4__slave ( .q(n208), .qb(n260), .d(NPC_reg_4__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n40), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_5__master ( .q(NPC_reg_5__m2s), .qb(), .d(N92), .sdi(n260),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_5__slave ( .q(n207), .qb(n259), .d(NPC_reg_5__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_6__master ( .q(NPC_reg_6__m2s), .qb(), .d(N93), .sdi(n259),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_6__slave ( .q(n206), .qb(n258), .d(NPC_reg_6__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 NPC_reg_7__master ( .q(NPC_reg_7__m2s), .qb(), .d(N94), .sdi(n258),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_4 NPC_reg_7__slave ( .q(NPC[7]), .qb(n26), .d(NPC_reg_7__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_8__master ( .q(NPC_reg_8__m2s), .qb(), .d(N95), .sdi(n26),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_8__slave ( .q(NPC[8]), .qb(n16), .d(NPC_reg_8__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_2 NPC_reg_9__master ( .q(NPC_reg_9__m2s), .qb(), .d(N96), .sdi(n16),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n36), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_8 NPC_reg_9__slave ( .q(NPC[9]), .qb(n22), .d(NPC_reg_9__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n36), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_0__master ( .q(PC_reg_0__m2s), .qb(), .d(n168), .sdi(n242),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_0__slave ( .q(PC[0]), .qb(n241), .d(PC_reg_0__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_10__master ( .q(PC_reg_10__m2s), .qb(), .d(n178), .sdi(n232),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_10__slave ( .q(PC[10]), .qb(n231), .d(PC_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_11__master ( .q(PC_reg_11__m2s), .qb(), .d(n179), .sdi(n231),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_11__slave ( .q(PC[11]), .qb(n230), .d(PC_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_12__master ( .q(PC_reg_12__m2s), .qb(), .d(n180), .sdi(n230),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_12__slave ( .q(PC[12]), .qb(n229), .d(PC_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_13__master ( .q(PC_reg_13__m2s), .qb(), .d(n181), .sdi(n229),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_13__slave ( .q(PC[13]), .qb(n228), .d(PC_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_14__master ( .q(PC_reg_14__m2s), .qb(), .d(n182), .sdi(n228),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_14__slave ( .q(PC[14]), .qb(n227), .d(PC_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_15__master ( .q(PC_reg_15__m2s), .qb(), .d(n183), .sdi(n227),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_15__slave ( .q(PC[15]), .qb(n226), .d(PC_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_16__master ( .q(PC_reg_16__m2s), .qb(), .d(n184), .sdi(n226),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n43), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_16__slave ( .q(PC[16]), .qb(n225), .d(PC_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n43), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_17__master ( .q(PC_reg_17__m2s), .qb(), .d(n185), .sdi(n225),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_17__slave ( .q(PC[17]), .qb(n224), .d(PC_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_18__master ( .q(PC_reg_18__m2s), .qb(), .d(n186), .sdi(n224),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_18__slave ( .q(PC[18]), .qb(n223), .d(PC_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_19__master ( .q(PC_reg_19__m2s), .qb(), .d(n187), .sdi(n223),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_19__slave ( .q(PC[19]), .qb(n222), .d(PC_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_1__master ( .q(PC_reg_1__m2s), .qb(), .d(n169), .sdi(n241),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_1__slave ( .q(PC[1]), .qb(n240), .d(PC_reg_1__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_20__master ( .q(PC_reg_20__m2s), .qb(), .d(n188), .sdi(n222),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_20__slave ( .q(PC[20]), .qb(n221), .d(PC_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_21__master ( .q(PC_reg_21__m2s), .qb(), .d(n189), .sdi(n221),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_21__slave ( .q(PC[21]), .qb(n92), .d(PC_reg_21__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_22__master ( .q(PC_reg_22__m2s), .qb(), .d(n190), .sdi(PC[21]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_22__slave ( .q(PC[22]), .qb(n93), .d(PC_reg_22__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_23__master ( .q(PC_reg_23__m2s), .qb(), .d(n191), .sdi(PC[22]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_23__slave ( .q(PC[23]), .qb(n94), .d(PC_reg_23__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_24__master ( .q(PC_reg_24__m2s), .qb(), .d(n192), .sdi(PC[23]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_24__slave ( .q(PC[24]), .qb(n95), .d(PC_reg_24__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_25__master ( .q(PC_reg_25__m2s), .qb(), .d(n193), .sdi(PC[24]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_25__slave ( .q(PC[25]), .qb(n96), .d(PC_reg_25__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_26__master ( .q(PC_reg_26__m2s), .qb(), .d(n194), .sdi(PC[25]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_26__slave ( .q(PC[26]), .qb(n97), .d(PC_reg_26__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_27__master ( .q(PC_reg_27__m2s), .qb(), .d(n195), .sdi(PC[26]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_27__slave ( .q(PC[27]), .qb(n98), .d(PC_reg_27__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_28__master ( .q(PC_reg_28__m2s), .qb(), .d(n196), .sdi(PC[27]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_28__slave ( .q(PC[28]), .qb(n99), .d(PC_reg_28__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_29__master ( .q(PC_reg_29__m2s), .qb(), .d(n197), .sdi(PC[28]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_29__slave ( .q(PC[29]), .qb(n100), .d(PC_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_2__master ( .q(PC_reg_2__m2s), .qb(), .d(n170), .sdi(n240),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_2__slave ( .q(PC[2]), .qb(n239), .d(PC_reg_2__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_30__master ( .q(PC_reg_30__m2s), .qb(), .d(n198), .sdi(PC[29]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_30__slave ( .q(PC[30]), .qb(n101), .d(PC_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_31__master ( .q(PC_reg_31__m2s), .qb(), .d(n199), .sdi(PC[30]),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_31__slave ( .q(PC[31]), .qb(n102), .d(PC_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_3__master ( .q(PC_reg_3__m2s), .qb(), .d(n171), .sdi(n239),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_3__slave ( .q(PC[3]), .qb(n238), .d(PC_reg_3__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_4__master ( .q(PC_reg_4__m2s), .qb(), .d(n172), .sdi(n238),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_4__slave ( .q(PC[4]), .qb(n237), .d(PC_reg_4__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_5__master ( .q(PC_reg_5__m2s), .qb(), .d(n173), .sdi(n237),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_5__slave ( .q(PC[5]), .qb(n236), .d(PC_reg_5__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_6__master ( .q(PC_reg_6__m2s), .qb(), .d(n174), .sdi(n236),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_6__slave ( .q(PC[6]), .qb(n235), .d(PC_reg_6__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_7__master ( .q(PC_reg_7__m2s), .qb(), .d(n175), .sdi(n235),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_7__slave ( .q(PC[7]), .qb(n234), .d(PC_reg_7__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_8__master ( .q(PC_reg_8__m2s), .qb(), .d(n176), .sdi(n234),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_8__slave ( .q(PC[8]), .qb(n233), .d(PC_reg_8__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 PC_reg_9__master ( .q(PC_reg_9__m2s), .qb(), .d(n177), .sdi(n233),
		.se(test_se), .g(Ctrl__Regs_1__en1), .rb(n39), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 PC_reg_9__slave ( .q(PC[9]), .qb(n232), .d(PC_reg_9__m2s), .g(Ctrl__Regs_1__en2),
		.rb(n39), .glob_g(global_g2), .sync_sel(sync_sel) );
	nand2_2 U10 ( .x(n48), .a(branch_address[22]), .b(branch_sig) );
	mux2_2 U100 ( .x(n163), .d0(IR_curr_27), .sl(n87), .d1(IR[27]) );
	mux2_2 U101 ( .x(n164), .d0(IR_curr_28), .sl(n87), .d1(IR[28]) );
	mux2_2 U102 ( .x(n165), .d0(IR_curr_29), .sl(n87), .d1(IR[29]) );
	buf_3 U103 ( .x(n42), .a(n91) );
	mux2_2 U104 ( .x(n166), .d0(IR_curr_30), .sl(n87), .d1(IR[30]) );
	buf_3 U105 ( .x(n41), .a(n91) );
	inv_2 U106 ( .x(n81), .a(counter[0]) );
	inv_2 U107 ( .x(n83), .a(counter[1]) );
	mux2_2 U108 ( .x(n168), .d0(PC[0]), .sl(n89), .d1(n218) );
	mux2_2 U109 ( .x(n169), .d0(PC[1]), .sl(n89), .d1(NPC[1]) );
	nand2i_2 U11 ( .x(n49), .a(n93), .b(N152) );
	mux2_2 U110 ( .x(n170), .d0(PC[2]), .sl(n89), .d1(n33) );
	mux2_2 U111 ( .x(n171), .d0(PC[3]), .sl(n90), .d1(n31) );
	buf_3 U112 ( .x(n43), .a(n91) );
	mux2_3 U113 ( .x(n186), .d0(PC[18]), .sl(n89), .d1(NPC[18]) );
	mux2_3 U114 ( .x(n187), .d0(PC[19]), .sl(n90), .d1(NPC[19]) );
	mux2_3 U115 ( .x(n188), .d0(PC[20]), .sl(n89), .d1(NPC[20]) );
	mux2_2 U116 ( .x(n189), .d0(PC[21]), .sl(n90), .d1(n214) );
	mux2_2 U117 ( .x(n190), .d0(PC[22]), .sl(n90), .d1(NPC[22]) );
	mux2_2 U118 ( .x(n191), .d0(PC[23]), .sl(n89), .d1(NPC[23]) );
	mux2_2 U119 ( .x(n192), .d0(PC[24]), .sl(n90), .d1(NPC[24]) );
	ao222_1 U12 ( .x(N150), .a(IR_previous_31), .b(N152), .c(IR_curr_31), .d(n4),
		.e(IR[31]), .f(n202) );
	mux2_3 U120 ( .x(n193), .d0(PC[25]), .sl(n89), .d1(NPC[25]) );
	mux2_2 U121 ( .x(n194), .d0(PC[26]), .sl(n89), .d1(NPC[26]) );
	mux2_2 U122 ( .x(n195), .d0(PC[27]), .sl(n90), .d1(NPC[27]) );
	mux2_2 U123 ( .x(n196), .d0(PC[28]), .sl(n90), .d1(NPC[28]) );
	mux2_2 U124 ( .x(n197), .d0(PC[29]), .sl(n89), .d1(NPC[29]) );
	mux2_2 U125 ( .x(n198), .d0(PC[30]), .sl(n89), .d1(NPC[30]) );
	buf_3 U126 ( .x(n39), .a(n91) );
	mux2_2 U127 ( .x(n199), .d0(PC[31]), .sl(n89), .d1(NPC[31]) );
	oai21_1 U128 ( .x(n200), .a(n90), .b(test_so1), .c(n88) );
	ao222_1 U129 ( .x(N119), .a(IR_previous_0), .b(n5), .c(IR_curr_0), .d(n4),
		.e(IR[0]), .f(n202) );
	ao222_1 U13 ( .x(N148), .a(IR_previous_29), .b(N152), .c(IR_curr_29), .d(n4),
		.e(IR[29]), .f(n202) );
	ao222_1 U130 ( .x(N120), .a(IR_previous_1), .b(n5), .c(IR_curr_1), .d(n4),
		.e(IR[1]), .f(n202) );
	ao222_1 U131 ( .x(N121), .a(IR_previous_2), .b(n5), .c(IR_curr_2), .d(n4),
		.e(IR[2]), .f(n202) );
	ao222_1 U132 ( .x(N122), .a(IR_previous_3), .b(n5), .c(IR_curr_3), .d(n4),
		.e(IR[3]), .f(n202) );
	ao222_1 U133 ( .x(N123), .a(IR_previous_4), .b(n5), .c(IR_curr_4), .d(n4),
		.e(IR[4]), .f(n202) );
	ao222_1 U134 ( .x(N124), .a(IR_previous_5), .b(n5), .c(IR_curr_5), .d(n4),
		.e(IR[5]), .f(n202) );
	ao222_1 U135 ( .x(N125), .a(IR_previous_6), .b(n5), .c(IR_curr_6), .d(n4),
		.e(IR[6]), .f(n202) );
	ao222_1 U136 ( .x(N127), .a(IR_previous_8), .b(n5), .c(IR_curr_8), .d(n4),
		.e(IR[8]), .f(n202) );
	ao222_1 U137 ( .x(N128), .a(IR_previous_9), .b(n5), .c(IR_curr_9), .d(n4),
		.e(IR[9]), .f(n202) );
	ao222_1 U138 ( .x(N129), .a(IR_previous_10), .b(n5), .c(IR_curr_10), .d(n4),
		.e(IR[10]), .f(n202) );
	ao222_1 U139 ( .x(N130), .a(IR_previous_11), .b(n5), .c(IR_curr_11), .d(n4),
		.e(IR[11]), .f(n202) );
	ao222_1 U14 ( .x(N88), .a(PC[1]), .b(n5), .c(branch_address[1]), .d(n6),
		.e(N18), .f(N215) );
	ao222_1 U140 ( .x(N131), .a(IR_previous_12), .b(n5), .c(IR_curr_12), .d(n4),
		.e(IR[12]), .f(n202) );
	ao222_1 U141 ( .x(N132), .a(IR_previous_13), .b(n5), .c(IR_curr_13), .d(n4),
		.e(IR[13]), .f(n202) );
	ao222_1 U142 ( .x(N133), .a(IR_previous_14), .b(n5), .c(IR_curr_14), .d(n4),
		.e(IR[14]), .f(n202) );
	ao222_1 U143 ( .x(N134), .a(IR_previous_15), .b(n5), .c(IR_curr_15), .d(n4),
		.e(IR[15]), .f(n202) );
	ao222_1 U144 ( .x(N135), .a(IR_previous_16), .b(n5), .c(IR_curr_16), .d(n4),
		.e(IR[16]), .f(n202) );
	ao222_1 U145 ( .x(N136), .a(IR_previous_17), .b(n5), .c(IR_curr_17), .d(n4),
		.e(IR[17]), .f(n202) );
	ao222_1 U146 ( .x(N137), .a(IR_previous_18), .b(n5), .c(IR_curr_18), .d(n4),
		.e(IR[18]), .f(n202) );
	ao222_1 U147 ( .x(N139), .a(IR_previous_20), .b(n5), .c(IR_curr_20), .d(n4),
		.e(IR[20]), .f(n202) );
	ao222_1 U148 ( .x(N140), .a(IR_previous_21), .b(n5), .c(IR_curr_21), .d(n4),
		.e(IR[21]), .f(n202) );
	ao222_1 U149 ( .x(N141), .a(IR_previous_22), .b(n5), .c(IR_curr_22), .d(n4),
		.e(IR[22]), .f(n202) );
	oai211_1 U15 ( .x(N108), .a(n201), .b(n44), .c(n45), .d(n46) );
	ao222_1 U150 ( .x(N142), .a(IR_previous_23), .b(n5), .c(IR_curr_23), .d(n4),
		.e(IR[23]), .f(n202) );
	ao222_1 U151 ( .x(N143), .a(IR_previous_24), .b(n5), .c(IR_curr_24), .d(n4),
		.e(IR[24]), .f(n202) );
	ao222_1 U152 ( .x(N144), .a(IR_previous_25), .b(n5), .c(IR_curr_25), .d(n4),
		.e(IR[25]), .f(n202) );
	ao222_1 U153 ( .x(N146), .a(IR_previous_27), .b(n5), .c(IR_curr_27), .d(n4),
		.e(IR[27]), .f(n202) );
	ao222_1 U154 ( .x(N147), .a(IR_previous_28), .b(n5), .c(IR_curr_28), .d(n4),
		.e(IR[28]), .f(n202) );
	buf_3 U155 ( .x(n37), .a(n91) );
	oai21_2 U156 ( .x(n202), .a(N50), .b(n201), .c(n203) );
	ao222_1 U157 ( .x(N149), .a(IR_previous_30), .b(n5), .c(IR_curr_30), .d(n4),
		.e(IR[30]), .f(n202) );
	nand2i_2 U158 ( .x(n61), .a(n97), .b(N152) );
	inv_2 U159 ( .x(n59), .a(N43) );
	inv_2 U16 ( .x(n44), .a(N38) );
	oai211_1 U160 ( .x(N113), .a(n201), .b(n59), .c(n60), .d(n61) );
	nand2i_2 U161 ( .x(n64), .a(n98), .b(N152) );
	nand2_2 U162 ( .x(n63), .a(branch_address[27]), .b(branch_sig) );
	inv_2 U163 ( .x(n62), .a(N44) );
	oai211_1 U164 ( .x(N114), .a(n201), .b(n62), .c(n63), .d(n64) );
	nand2i_2 U165 ( .x(n67), .a(n99), .b(N152) );
	nand2_2 U166 ( .x(n66), .a(branch_address[28]), .b(branch_sig) );
	inv_2 U167 ( .x(n65), .a(N45) );
	oai211_1 U168 ( .x(N115), .a(n201), .b(n65), .c(n66), .d(n67) );
	inv_2 U169 ( .x(n86), .a(n69) );
	nand2_2 U17 ( .x(n45), .a(branch_address[21]), .b(branch_sig) );
	nor2i_1 U170 ( .x(n70), .a(n68), .b(n86) );
	nand2i_2 U171 ( .x(n69), .a(n100), .b(N152) );
	nand2_2 U172 ( .x(n68), .a(branch_address[29]), .b(branch_sig) );
	inv_2 U173 ( .x(n85), .a(n78) );
	nor2i_1 U174 ( .x(n79), .a(n77), .b(n85) );
	nand2_2 U175 ( .x(n77), .a(branch_address[30]), .b(branch_sig) );
	inv_2 U176 ( .x(n89), .a(n201) );
	inv_2 U177 ( .x(n90), .a(n201) );
	inv_5 U178 ( .x(n76), .a(N48) );
	inv_2 U179 ( .x(n84), .a(n74) );
	nand2i_2 U18 ( .x(n46), .a(n92), .b(N152) );
	nor2i_1 U180 ( .x(n75), .a(n73), .b(n84) );
	nand2_2 U181 ( .x(n73), .a(branch_address[31]), .b(branch_sig) );
	aoi23_1 U182 ( .x(N118), .a(n75), .b(n76), .c(n73), .d(n201), .e(n74) );
	buf_14 U183 ( .x(NPC[4]), .a(n208) );
	inv_2 U184 ( .x(n82), .a(stall) );
	and2_3 U185 ( .x(n4), .a(N50), .b(N215) );
	buf_3 U186 ( .x(n40), .a(n91) );
	buf_3 U187 ( .x(n38), .a(n91) );
	inv_5 U188 ( .x(N152), .a(n88) );
	inv_2 U189 ( .x(n5), .a(n88) );
	ao222_1 U19 ( .x(N138), .a(IR_previous_19), .b(N152), .c(IR_curr_19), .d(n4),
		.e(IR[19]), .f(n202) );
	nand2i_2 U190 ( .x(n88), .a(branch_sig), .b(n72) );
	ao222_1 U191 ( .x(N104), .a(PC[17]), .b(N152), .c(branch_address[17]),
		.d(n6), .e(N34), .f(N215) );
	ao222_1 U192 ( .x(N98), .a(PC[11]), .b(N152), .c(branch_address[11]), .d(branch_sig),
		.e(N28), .f(N215) );
	inv_2 U193 ( .x(n6), .a(n203) );
	inv_2 U194 ( .x(n203), .a(branch_sig) );
	inv_2 U195 ( .x(n8), .a(n72) );
	inv_2 U196 ( .x(n7), .a(n72) );
	inv_2 U197 ( .x(n87), .a(n72) );
	nand3_1 U198 ( .x(n72), .a(n81), .b(n82), .c(n83) );
	buf_14 U199 ( .x(NPC[15]), .a(n204) );
	oai211_1 U20 ( .x(N112), .a(n201), .b(n56), .c(n57), .d(n58) );
	ao222_1 U201 ( .x(N92), .a(PC[5]), .b(N152), .c(branch_address[5]), .d(branch_sig),
		.e(N22), .f(N215) );
	ao222_1 U202 ( .x(N101), .a(PC[14]), .b(N152), .c(branch_address[14]),
		.d(branch_sig), .e(N31), .f(N215) );
	inv_2 U203 ( .x(n11), .a(n10) );
	buf_10 U204 ( .x(NPC[11]), .a(n205) );
	inv_2 U205 ( .x(n13), .a(n12) );
	inv_2 U206 ( .x(n15), .a(n14) );
	mux2_1 U207 ( .x(n184), .d0(PC[16]), .sl(n90), .d1(NPC[16]) );
	ao222_1 U208 ( .x(N87), .a(PC[0]), .b(N152), .c(branch_address[0]), .d(branch_sig),
		.e(N17), .f(N215) );
	ao222_1 U209 ( .x(N91), .a(PC[4]), .b(N152), .c(branch_address[4]), .d(branch_sig),
		.e(N21), .f(N215) );
	inv_2 U21 ( .x(n56), .a(N42) );
	ao222_1 U210 ( .x(N97), .a(PC[10]), .b(N152), .c(branch_address[10]), .d(branch_sig),
		.e(N27), .f(N215) );
	ao222_1 U211 ( .x(N93), .a(PC[6]), .b(N152), .c(branch_address[6]), .d(branch_sig),
		.e(N23), .f(N215) );
	nand2_2 U212 ( .x(n60), .a(branch_address[26]), .b(branch_sig) );
	inv_2 U214 ( .x(n17), .a(n16) );
	mux2_1 U215 ( .x(n183), .d0(PC[15]), .sl(n89), .d1(NPC[15]) );
	mux2_1 U216 ( .x(n185), .d0(PC[17]), .sl(n90), .d1(n11) );
	mux2_1 U217 ( .x(n176), .d0(PC[8]), .sl(n89), .d1(n17) );
	inv_2 U218 ( .x(n23), .a(n22) );
	mux2_1 U219 ( .x(n174), .d0(PC[6]), .sl(n89), .d1(n211) );
	nand2_2 U22 ( .x(n57), .a(branch_address[25]), .b(branch_sig) );
	inv_2 U220 ( .x(n25), .a(n24) );
	inv_2 U221 ( .x(n27), .a(n26) );
	mux2_1 U222 ( .x(n181), .d0(PC[13]), .sl(n90), .d1(n15) );
	mux2_1 U223 ( .x(n172), .d0(PC[4]), .sl(n90), .d1(NPC[4]) );
	mux2_1 U224 ( .x(n182), .d0(PC[14]), .sl(n89), .d1(n13) );
	ao222_1 U225 ( .x(N90), .a(PC[3]), .b(N152), .c(branch_address[3]), .d(branch_sig),
		.e(N20), .f(N215) );
	mux2_1 U226 ( .x(n178), .d0(PC[10]), .sl(n89), .d1(n25) );
	inv_2 U227 ( .x(n29), .a(n28) );
	inv_2 U228 ( .x(n31), .a(n30) );
	inv_2 U229 ( .x(n33), .a(n32) );
	nand2i_2 U23 ( .x(n58), .a(n96), .b(N152) );
	mux2_1 U230 ( .x(n179), .d0(PC[11]), .sl(n90), .d1(NPC[11]) );
	mux2_1 U231 ( .x(n177), .d0(PC[9]), .sl(n89), .d1(n23) );
	mux2_1 U232 ( .x(n175), .d0(PC[7]), .sl(n90), .d1(n27) );
	mux2_1 U233 ( .x(n180), .d0(PC[12]), .sl(n89), .d1(n29) );
	buf_16 U234 ( .x(NPC[3]), .a(n209) );
	buf_16 U235 ( .x(NPC[2]), .a(n210) );
	mux2_1 U236 ( .x(n173), .d0(PC[5]), .sl(n90), .d1(n212) );
	inv_6 U237 ( .x(n71), .a(N46) );
	inv_6 U238 ( .x(n80), .a(N47) );
	nand2i_4 U239 ( .x(n74), .a(n102), .b(N152) );
	ao222_1 U24 ( .x(N126), .a(IR_previous_7), .b(N152), .c(IR_curr_7), .d(n4),
		.e(IR[7]), .f(n202) );
	nand2i_4 U240 ( .x(n78), .a(n101), .b(N152) );
	nand2i_6 U241 ( .x(n201), .a(branch_sig), .b(n7) );
	aoi23_4 U242 ( .x(N116), .a(n70), .b(n71), .c(n68), .d(n201), .e(n69) );
	aoi23_4 U243 ( .x(N117), .a(n79), .b(n80), .c(n77), .d(n201), .e(n78) );
	mux2_4 U244 ( .x(n167), .d0(IR_curr_31), .sl(n87), .d1(IR[31]) );
	inv_2 U245 ( .x(n91), .a(reset) );
	ao222_5 U247 ( .x(N99), .a(N152), .b(PC[12]), .c(branch_sig), .d(branch_address[12]),
		.e(N29), .f(N215) );
	inv_2 U248 ( .x(n211), .a(n258) );
	buf_10 U249 ( .x(NPC[6]), .a(n206) );
	ao222_2 U25 ( .x(N107), .a(PC[20]), .b(n5), .c(branch_address[20]), .d(n6),
		.e(N37), .f(N215) );
	inv_2 U250 ( .x(n212), .a(n259) );
	buf_10 U251 ( .x(NPC[5]), .a(n207) );
	inv_0 U252 ( .x(n213), .a(NPC[21]) );
	inv_2 U253 ( .x(n214), .a(n213) );
	inv_5 U254 ( .x(n215), .a(n360) );
	inv_10 U255 ( .x(NPC[14]), .a(n215) );
	ao222_1 U256 ( .x(N103), .a(PC[16]), .b(n5), .c(branch_address[16]), .d(branch_sig),
		.e(N33), .f(N215) );
	inv_0 U257 ( .x(n217), .a(NPC[0]) );
	inv_2 U258 ( .x(n218), .a(n217) );
	ao222_1 U259 ( .x(N100), .a(PC[13]), .b(N152), .c(branch_address[13]),
		.d(branch_sig), .e(N30), .f(N215) );
	oai211_1 U26 ( .x(N110), .a(n201), .b(n50), .c(n51), .d(n52) );
	ao222_1 U260 ( .x(N106), .a(PC[19]), .b(N152), .c(branch_address[19]),
		.d(branch_sig), .e(N36), .f(N215) );
	inv_5 U27 ( .x(n50), .a(N40) );
	nand2_2 U28 ( .x(n51), .a(branch_address[23]), .b(branch_sig) );
	nand2i_2 U29 ( .x(n52), .a(n94), .b(N152) );
	oai211_1 U3 ( .x(N111), .a(n201), .b(n53), .c(n54), .d(n55) );
	inv_2 U30 ( .x(N215), .a(n201) );
	ao222_1 U31 ( .x(N105), .a(PC[18]), .b(N152), .c(branch_address[18]), .d(branch_sig),
		.e(N35), .f(N215) );
	ao222_1 U32 ( .x(N145), .a(IR_previous_26), .b(N152), .c(IR_curr_26), .d(n4),
		.e(IR[26]), .f(n202) );
	ao222_1 U33 ( .x(N102), .a(PC[15]), .b(n5), .c(branch_address[15]), .d(branch_sig),
		.e(N32), .f(N215) );
	ao222_4 U36 ( .x(N94), .a(PC[7]), .b(N152), .c(branch_address[7]), .d(branch_sig),
		.e(N24), .f(N215) );
	ao222_4 U37 ( .x(N96), .a(PC[9]), .b(n5), .c(branch_address[9]), .d(branch_sig),
		.e(N26), .f(N215) );
	ao222_1 U38 ( .x(N95), .a(PC[8]), .b(N152), .c(branch_address[8]), .d(branch_sig),
		.e(N25), .f(N215) );
	buf_3 U39 ( .x(n36), .a(n91) );
	ao222_1 U40 ( .x(N89), .a(PC[2]), .b(N152), .c(branch_address[2]), .d(branch_sig),
		.e(N19), .f(N215) );
	mux2_2 U41 ( .x(n104), .d0(IR_previous_0), .sl(n8), .d1(IR_latched[0]) );
	mux2_2 U42 ( .x(n105), .d0(IR_previous_1), .sl(n8), .d1(IR_latched[1]) );
	mux2_2 U43 ( .x(n106), .d0(IR_previous_2), .sl(n8), .d1(IR_latched[2]) );
	mux2_2 U44 ( .x(n107), .d0(IR_previous_3), .sl(n87), .d1(IR_latched[3]) );
	mux2_2 U45 ( .x(n108), .d0(IR_previous_4), .sl(n8), .d1(IR_latched[4]) );
	mux2_2 U46 ( .x(n109), .d0(IR_previous_5), .sl(n87), .d1(IR_latched[5]) );
	mux2_2 U47 ( .x(n110), .d0(IR_previous_6), .sl(n8), .d1(IR_latched[6]) );
	mux2_2 U48 ( .x(n111), .d0(IR_previous_7), .sl(n87), .d1(IR_latched[7]) );
	mux2_2 U49 ( .x(n112), .d0(IR_previous_8), .sl(n87), .d1(IR_latched[8]) );
	inv_2 U5 ( .x(n53), .a(N41) );
	mux2_2 U50 ( .x(n113), .d0(IR_previous_9), .sl(n87), .d1(IR_latched[9]) );
	mux2_2 U51 ( .x(n114), .d0(IR_previous_10), .sl(n8), .d1(IR_latched[10]) );
	mux2_2 U52 ( .x(n115), .d0(IR_previous_11), .sl(n8), .d1(IR_latched[11]) );
	mux2_2 U53 ( .x(n116), .d0(IR_previous_12), .sl(n8), .d1(IR_latched[12]) );
	mux2_2 U54 ( .x(n117), .d0(IR_previous_13), .sl(n8), .d1(IR_latched[13]) );
	mux2_2 U55 ( .x(n118), .d0(IR_previous_14), .sl(n8), .d1(IR_latched[14]) );
	mux2_2 U56 ( .x(n119), .d0(IR_previous_15), .sl(n87), .d1(IR_latched[15]) );
	mux2_2 U57 ( .x(n120), .d0(IR_previous_16), .sl(n8), .d1(IR_latched[16]) );
	mux2_2 U58 ( .x(n121), .d0(IR_previous_17), .sl(n87), .d1(IR_latched[17]) );
	mux2_2 U59 ( .x(n122), .d0(IR_previous_18), .sl(n8), .d1(IR_latched[18]) );
	nand2_2 U6 ( .x(n54), .a(branch_address[24]), .b(branch_sig) );
	mux2_2 U60 ( .x(n123), .d0(IR_previous_19), .sl(n87), .d1(IR_latched[19]) );
	mux2_2 U61 ( .x(n124), .d0(IR_previous_20), .sl(n87), .d1(IR_latched[20]) );
	mux2_2 U62 ( .x(n125), .d0(IR_previous_21), .sl(n8), .d1(IR_latched[21]) );
	mux2_2 U63 ( .x(n126), .d0(IR_previous_22), .sl(n87), .d1(IR_latched[22]) );
	mux2_2 U64 ( .x(n127), .d0(IR_previous_23), .sl(n8), .d1(IR_latched[23]) );
	mux2_2 U65 ( .x(n128), .d0(IR_previous_24), .sl(n87), .d1(IR_latched[24]) );
	mux2_2 U66 ( .x(n129), .d0(IR_previous_25), .sl(n8), .d1(IR_latched[25]) );
	mux2_2 U67 ( .x(n130), .d0(IR_previous_26), .sl(n87), .d1(IR_latched[26]) );
	mux2_2 U68 ( .x(n131), .d0(IR_previous_27), .sl(n8), .d1(IR_latched[27]) );
	mux2_2 U69 ( .x(n132), .d0(IR_previous_28), .sl(n87), .d1(IR_latched[28]) );
	nand2i_2 U7 ( .x(n55), .a(n95), .b(N152) );
	mux2_2 U70 ( .x(n133), .d0(IR_previous_29), .sl(n8), .d1(IR_latched[29]) );
	mux2_2 U71 ( .x(n134), .d0(IR_previous_30), .sl(n8), .d1(IR_latched[30]) );
	mux2_2 U72 ( .x(n135), .d0(IR_previous_31), .sl(n87), .d1(IR_latched[31]) );
	mux2_2 U73 ( .x(n136), .d0(IR_curr_0), .sl(n8), .d1(IR[0]) );
	mux2_2 U74 ( .x(n137), .d0(IR_curr_1), .sl(n8), .d1(IR[1]) );
	mux2_2 U75 ( .x(n138), .d0(IR_curr_2), .sl(n87), .d1(IR[2]) );
	mux2_2 U76 ( .x(n139), .d0(IR_curr_3), .sl(n87), .d1(IR[3]) );
	mux2_2 U77 ( .x(n140), .d0(IR_curr_4), .sl(n87), .d1(IR[4]) );
	mux2_2 U78 ( .x(n141), .d0(IR_curr_5), .sl(n87), .d1(IR[5]) );
	mux2_2 U79 ( .x(n142), .d0(IR_curr_6), .sl(n87), .d1(IR[6]) );
	oai211_1 U8 ( .x(N109), .a(n201), .b(n47), .c(n48), .d(n49) );
	mux2_2 U80 ( .x(n143), .d0(IR_curr_7), .sl(n87), .d1(IR[7]) );
	mux2_2 U81 ( .x(n144), .d0(IR_curr_8), .sl(n87), .d1(IR[8]) );
	mux2_2 U82 ( .x(n145), .d0(IR_curr_9), .sl(n87), .d1(IR[9]) );
	mux2_2 U83 ( .x(n146), .d0(IR_curr_10), .sl(n8), .d1(IR[10]) );
	mux2_2 U84 ( .x(n147), .d0(IR_curr_11), .sl(n8), .d1(IR[11]) );
	mux2_2 U85 ( .x(n148), .d0(IR_curr_12), .sl(n8), .d1(IR[12]) );
	mux2_2 U86 ( .x(n149), .d0(IR_curr_13), .sl(n8), .d1(IR[13]) );
	mux2_2 U87 ( .x(n150), .d0(IR_curr_14), .sl(n8), .d1(IR[14]) );
	mux2_2 U88 ( .x(n151), .d0(IR_curr_15), .sl(n8), .d1(IR[15]) );
	mux2_2 U89 ( .x(n152), .d0(IR_curr_16), .sl(n8), .d1(IR[16]) );
	inv_2 U9 ( .x(n47), .a(N39) );
	mux2_2 U90 ( .x(n153), .d0(IR_curr_17), .sl(n8), .d1(IR[17]) );
	mux2_2 U91 ( .x(n154), .d0(IR_curr_18), .sl(n8), .d1(IR[18]) );
	mux2_2 U92 ( .x(n155), .d0(IR_curr_19), .sl(n87), .d1(IR[19]) );
	mux2_2 U93 ( .x(n156), .d0(IR_curr_20), .sl(n87), .d1(IR[20]) );
	mux2_2 U94 ( .x(n157), .d0(IR_curr_21), .sl(n87), .d1(IR[21]) );
	mux2_2 U95 ( .x(n158), .d0(IR_curr_22), .sl(n8), .d1(IR[22]) );
	mux2_2 U96 ( .x(n159), .d0(IR_curr_23), .sl(n8), .d1(IR[23]) );
	mux2_2 U97 ( .x(n160), .d0(IR_curr_24), .sl(n8), .d1(IR[24]) );
	mux2_2 U98 ( .x(n161), .d0(IR_curr_25), .sl(n87), .d1(IR[25]) );
	mux2_2 U99 ( .x(n162), .d0(IR_curr_26), .sl(n87), .d1(IR[26]) );
	IF_DW01_add_32_0_test_1 add_100 ( .A({ NPC[31], NPC[30], NPC[29], NPC[28],
		NPC[27], NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], n214, NPC[20],
		NPC[19], NPC[18], n11, NPC[16], NPC[15], n13, n15, n29, NPC[11], n25,
		n23, n17, n27, n211, n212, NPC[4], n31, n33, NPC[1], n218}), .B({ 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0,
		1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM({ N48, N47,
		N46, N45, N44, N43, N42, N41, N40, N39, N38, N37, N36, N35, N34, N33,
		N32, N31, N30, N29, N28, N27, N26, N25, N24, N23, N22, N21, N20, N19,
		N18, N17}), .CO() );
	smlatnr_1 stalled_reg__master ( .q(stalled_reg__m2s), .qb(), .d(n200),
		.sdi(PC[31]), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n38), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 stalled_reg__slave ( .q(N50), .qb(test_so1), .d(stalled_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n38), .glob_g(global_g2), .sync_sel(sync_sel) );

endmodule


module MEM_test_1_desync (  reg_write_MEM, mem_to_reg_EX, reset, ALU_result,
	reg_write_EX, mem_to_reg_MEM, reg_out_B_EX, reg_out_B_MEM, DM_read_data,
	RF_data_in, test_si, test_so, test_se, sync_sel, global_g1, global_g2,
	Ctrl__Regs_1__en1, Ctrl__Regs_1__en2 );

input  mem_to_reg_EX, reset, reg_write_EX, test_si, test_se, sync_sel, global_g1,
	global_g2, Ctrl__Regs_1__en1, Ctrl__Regs_1__en2;
input [31:0] ALU_result, reg_out_B_EX, DM_read_data;
output  reg_write_MEM, mem_to_reg_MEM, test_so;
output [31:0] reg_out_B_MEM, RF_data_in;

wire RF_data_in_reg_0__m2s, RF_data_in_reg_10__m2s, RF_data_in_reg_11__m2s,
	RF_data_in_reg_12__m2s, RF_data_in_reg_13__m2s, RF_data_in_reg_14__m2s,
	RF_data_in_reg_15__m2s, RF_data_in_reg_16__m2s, RF_data_in_reg_17__m2s,
	RF_data_in_reg_18__m2s, RF_data_in_reg_19__m2s, RF_data_in_reg_1__m2s,
	RF_data_in_reg_20__m2s, RF_data_in_reg_21__m2s, RF_data_in_reg_22__m2s,
	RF_data_in_reg_23__m2s, RF_data_in_reg_24__m2s, RF_data_in_reg_25__m2s,
	RF_data_in_reg_26__m2s, RF_data_in_reg_27__m2s, RF_data_in_reg_28__m2s,
	RF_data_in_reg_29__m2s, RF_data_in_reg_2__m2s, RF_data_in_reg_30__m2s,
	RF_data_in_reg_31__m2s, RF_data_in_reg_3__m2s, RF_data_in_reg_4__m2s,
	RF_data_in_reg_5__m2s, RF_data_in_reg_6__m2s, RF_data_in_reg_7__m2s, RF_data_in_reg_8__m2s,
	RF_data_in_reg_9__m2s, mem_to_reg_MEM_reg__m2s, n11, n12, n13, n14, n15,
	n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
	n3, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n4, n40, n41, n42,
	n43, n44, n45, n46, n47, n48, n49, n5, n50, n51, n52, n53, n54, n55, n56,
	n57, n58, n59, n6, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
	n71, n72, n73, n74, n75, reg_out_B_MEM_reg_0__m2s, reg_out_B_MEM_reg_10__m2s,
	reg_out_B_MEM_reg_11__m2s, reg_out_B_MEM_reg_12__m2s, reg_out_B_MEM_reg_13__m2s,
	reg_out_B_MEM_reg_14__m2s, reg_out_B_MEM_reg_15__m2s, reg_out_B_MEM_reg_16__m2s,
	reg_out_B_MEM_reg_17__m2s, reg_out_B_MEM_reg_18__m2s, reg_out_B_MEM_reg_19__m2s,
	reg_out_B_MEM_reg_1__m2s, reg_out_B_MEM_reg_20__m2s, reg_out_B_MEM_reg_21__m2s,
	reg_out_B_MEM_reg_22__m2s, reg_out_B_MEM_reg_23__m2s, reg_out_B_MEM_reg_24__m2s,
	reg_out_B_MEM_reg_25__m2s, reg_out_B_MEM_reg_26__m2s, reg_out_B_MEM_reg_27__m2s,
	reg_out_B_MEM_reg_28__m2s, reg_out_B_MEM_reg_29__m2s, reg_out_B_MEM_reg_2__m2s,
	reg_out_B_MEM_reg_30__m2s, reg_out_B_MEM_reg_31__m2s, reg_out_B_MEM_reg_3__m2s,
	reg_out_B_MEM_reg_4__m2s, reg_out_B_MEM_reg_5__m2s, reg_out_B_MEM_reg_6__m2s,
	reg_out_B_MEM_reg_7__m2s, reg_out_B_MEM_reg_8__m2s, reg_out_B_MEM_reg_9__m2s,
	reg_write_MEM_reg__m2s;


	smlatnr_1 RF_data_in_reg_0__master ( .q(RF_data_in_reg_0__m2s), .qb(),
		.d(n15), .sdi(test_si), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4),
		.glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 RF_data_in_reg_0__slave ( .q(RF_data_in[0]), .qb(n16), .d(RF_data_in_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_10__master ( .q(RF_data_in_reg_10__m2s), .qb(),
		.d(n69), .sdi(n18), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_10__slave ( .q(RF_data_in[10]), .qb(n70), .d(RF_data_in_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_11__master ( .q(RF_data_in_reg_11__m2s), .qb(),
		.d(n43), .sdi(n70), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_11__slave ( .q(RF_data_in[11]), .qb(n44), .d(RF_data_in_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_12__master ( .q(RF_data_in_reg_12__m2s), .qb(),
		.d(n67), .sdi(n44), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_12__slave ( .q(RF_data_in[12]), .qb(n68), .d(RF_data_in_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_13__master ( .q(RF_data_in_reg_13__m2s), .qb(),
		.d(n65), .sdi(n68), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_13__slave ( .q(RF_data_in[13]), .qb(n66), .d(RF_data_in_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_14__master ( .q(RF_data_in_reg_14__m2s), .qb(),
		.d(n11), .sdi(n66), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_14__slave ( .q(RF_data_in[14]), .qb(n12), .d(RF_data_in_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_15__master ( .q(RF_data_in_reg_15__m2s), .qb(),
		.d(n63), .sdi(n12), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_15__slave ( .q(RF_data_in[15]), .qb(n64), .d(RF_data_in_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_16__master ( .q(RF_data_in_reg_16__m2s), .qb(),
		.d(n61), .sdi(n64), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_16__slave ( .q(RF_data_in[16]), .qb(n62), .d(RF_data_in_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_17__master ( .q(RF_data_in_reg_17__m2s), .qb(),
		.d(n59), .sdi(n62), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_17__slave ( .q(RF_data_in[17]), .qb(n60), .d(RF_data_in_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_18__master ( .q(RF_data_in_reg_18__m2s), .qb(),
		.d(n57), .sdi(n60), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_18__slave ( .q(RF_data_in[18]), .qb(n58), .d(RF_data_in_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_19__master ( .q(RF_data_in_reg_19__m2s), .qb(),
		.d(n35), .sdi(n58), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_19__slave ( .q(RF_data_in[19]), .qb(n36), .d(RF_data_in_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_1__master ( .q(RF_data_in_reg_1__m2s), .qb(),
		.d(n13), .sdi(n16), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 RF_data_in_reg_1__slave ( .q(RF_data_in[1]), .qb(n14), .d(RF_data_in_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_20__master ( .q(RF_data_in_reg_20__m2s), .qb(),
		.d(n55), .sdi(n36), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_20__slave ( .q(RF_data_in[20]), .qb(n56), .d(RF_data_in_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_21__master ( .q(RF_data_in_reg_21__m2s), .qb(),
		.d(n53), .sdi(n56), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_21__slave ( .q(RF_data_in[21]), .qb(n54), .d(RF_data_in_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_22__master ( .q(RF_data_in_reg_22__m2s), .qb(),
		.d(n33), .sdi(n54), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_22__slave ( .q(RF_data_in[22]), .qb(n34), .d(RF_data_in_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_23__master ( .q(RF_data_in_reg_23__m2s), .qb(),
		.d(n51), .sdi(n34), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_23__slave ( .q(RF_data_in[23]), .qb(n52), .d(RF_data_in_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_24__master ( .q(RF_data_in_reg_24__m2s), .qb(),
		.d(n49), .sdi(n52), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_24__slave ( .q(RF_data_in[24]), .qb(n50), .d(RF_data_in_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_25__master ( .q(RF_data_in_reg_25__m2s), .qb(),
		.d(n47), .sdi(n50), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_25__slave ( .q(RF_data_in[25]), .qb(n48), .d(RF_data_in_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_26__master ( .q(RF_data_in_reg_26__m2s), .qb(),
		.d(n21), .sdi(n48), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_26__slave ( .q(RF_data_in[26]), .qb(n22), .d(RF_data_in_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_27__master ( .q(RF_data_in_reg_27__m2s), .qb(),
		.d(n31), .sdi(n22), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_27__slave ( .q(RF_data_in[27]), .qb(n32), .d(RF_data_in_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_28__master ( .q(RF_data_in_reg_28__m2s), .qb(),
		.d(n45), .sdi(n32), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_28__slave ( .q(RF_data_in[28]), .qb(n46), .d(RF_data_in_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_29__master ( .q(RF_data_in_reg_29__m2s), .qb(),
		.d(n29), .sdi(n46), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_29__slave ( .q(RF_data_in[29]), .qb(n30), .d(RF_data_in_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_2__master ( .q(RF_data_in_reg_2__m2s), .qb(),
		.d(n39), .sdi(n14), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 RF_data_in_reg_2__slave ( .q(RF_data_in[2]), .qb(n40), .d(RF_data_in_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_30__master ( .q(RF_data_in_reg_30__m2s), .qb(),
		.d(n25), .sdi(n30), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_30__slave ( .q(RF_data_in[30]), .qb(n26), .d(RF_data_in_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_31__master ( .q(RF_data_in_reg_31__m2s), .qb(),
		.d(n23), .sdi(n26), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_31__slave ( .q(RF_data_in[31]), .qb(n24), .d(RF_data_in_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_3__master ( .q(RF_data_in_reg_3__m2s), .qb(),
		.d(n41), .sdi(n40), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 RF_data_in_reg_3__slave ( .q(RF_data_in[3]), .qb(n42), .d(RF_data_in_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_4__master ( .q(RF_data_in_reg_4__m2s), .qb(),
		.d(n73), .sdi(n42), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 RF_data_in_reg_4__slave ( .q(RF_data_in[4]), .qb(n74), .d(RF_data_in_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_5__master ( .q(RF_data_in_reg_5__m2s), .qb(),
		.d(n71), .sdi(n74), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 RF_data_in_reg_5__slave ( .q(RF_data_in[5]), .qb(n72), .d(RF_data_in_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_6__master ( .q(RF_data_in_reg_6__m2s), .qb(),
		.d(n37), .sdi(n72), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n4), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 RF_data_in_reg_6__slave ( .q(RF_data_in[6]), .qb(n38), .d(RF_data_in_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_7__master ( .q(RF_data_in_reg_7__m2s), .qb(),
		.d(n19), .sdi(n38), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_4 RF_data_in_reg_7__slave ( .q(n75), .qb(n20), .d(RF_data_in_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_8__master ( .q(RF_data_in_reg_8__m2s), .qb(),
		.d(n27), .sdi(n20), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n6), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_8__slave ( .q(RF_data_in[8]), .qb(n28), .d(RF_data_in_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 RF_data_in_reg_9__master ( .q(RF_data_in_reg_9__m2s), .qb(),
		.d(n17), .sdi(n28), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_1 RF_data_in_reg_9__slave ( .q(RF_data_in[9]), .qb(n18), .d(RF_data_in_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	mux2_1 U10 ( .x(n23), .d0(ALU_result[31]), .sl(mem_to_reg_EX), .d1(DM_read_data[31]) );
	mux2_1 U11 ( .x(n25), .d0(ALU_result[30]), .sl(mem_to_reg_EX), .d1(DM_read_data[30]) );
	mux2_1 U12 ( .x(n27), .d0(ALU_result[8]), .sl(mem_to_reg_EX), .d1(DM_read_data[8]) );
	mux2_1 U13 ( .x(n29), .d0(ALU_result[29]), .sl(mem_to_reg_EX), .d1(DM_read_data[29]) );
	mux2_1 U14 ( .x(n31), .d0(ALU_result[27]), .sl(mem_to_reg_EX), .d1(DM_read_data[27]) );
	mux2_1 U15 ( .x(n33), .d0(ALU_result[22]), .sl(mem_to_reg_EX), .d1(DM_read_data[22]) );
	mux2_1 U16 ( .x(n35), .d0(ALU_result[19]), .sl(mem_to_reg_EX), .d1(DM_read_data[19]) );
	mux2_1 U17 ( .x(n37), .d0(ALU_result[6]), .sl(mem_to_reg_EX), .d1(DM_read_data[6]) );
	mux2_1 U18 ( .x(n39), .d0(ALU_result[2]), .sl(mem_to_reg_EX), .d1(DM_read_data[2]) );
	mux2_1 U19 ( .x(n41), .d0(ALU_result[3]), .sl(mem_to_reg_EX), .d1(DM_read_data[3]) );
	mux2_1 U20 ( .x(n43), .d0(ALU_result[11]), .sl(mem_to_reg_EX), .d1(DM_read_data[11]) );
	mux2_1 U21 ( .x(n45), .d0(ALU_result[28]), .sl(mem_to_reg_EX), .d1(DM_read_data[28]) );
	mux2_1 U22 ( .x(n47), .d0(ALU_result[25]), .sl(mem_to_reg_EX), .d1(DM_read_data[25]) );
	mux2_1 U23 ( .x(n49), .d0(ALU_result[24]), .sl(mem_to_reg_EX), .d1(DM_read_data[24]) );
	mux2_1 U24 ( .x(n51), .d0(ALU_result[23]), .sl(mem_to_reg_EX), .d1(DM_read_data[23]) );
	mux2_1 U25 ( .x(n53), .d0(ALU_result[21]), .sl(mem_to_reg_EX), .d1(DM_read_data[21]) );
	mux2_1 U26 ( .x(n55), .d0(ALU_result[20]), .sl(mem_to_reg_EX), .d1(DM_read_data[20]) );
	mux2_1 U27 ( .x(n57), .d0(ALU_result[18]), .sl(mem_to_reg_EX), .d1(DM_read_data[18]) );
	mux2_1 U28 ( .x(n59), .d0(ALU_result[17]), .sl(mem_to_reg_EX), .d1(DM_read_data[17]) );
	mux2_1 U29 ( .x(n61), .d0(ALU_result[16]), .sl(mem_to_reg_EX), .d1(DM_read_data[16]) );
	buf_3 U3 ( .x(n3), .a(mem_to_reg_EX) );
	mux2_1 U30 ( .x(n63), .d0(ALU_result[15]), .sl(mem_to_reg_EX), .d1(DM_read_data[15]) );
	mux2_1 U31 ( .x(n65), .d0(ALU_result[13]), .sl(mem_to_reg_EX), .d1(DM_read_data[13]) );
	mux2_1 U32 ( .x(n67), .d0(ALU_result[12]), .sl(mem_to_reg_EX), .d1(DM_read_data[12]) );
	mux2_1 U33 ( .x(n69), .d0(ALU_result[10]), .sl(mem_to_reg_EX), .d1(DM_read_data[10]) );
	mux2_1 U34 ( .x(n71), .d0(ALU_result[5]), .sl(mem_to_reg_EX), .d1(DM_read_data[5]) );
	mux2_1 U35 ( .x(n73), .d0(ALU_result[4]), .sl(n3), .d1(DM_read_data[4]) );
	inv_2 U4 ( .x(n5), .a(reset) );
	inv_2 U5 ( .x(n4), .a(reset) );
	inv_2 U6 ( .x(n6), .a(reset) );
	buf_16 U7 ( .x(RF_data_in[7]), .a(n75) );
	mux2_1 U8 ( .x(n19), .d0(ALU_result[7]), .sl(mem_to_reg_EX), .d1(DM_read_data[7]) );
	mux2_1 U9 ( .x(n21), .d0(ALU_result[26]), .sl(mem_to_reg_EX), .d1(DM_read_data[26]) );
	mux2_1 _RF_data_in_reg_0_U4 ( .x(n15), .d0(ALU_result[0]), .sl(mem_to_reg_EX),
		.d1(DM_read_data[0]) );
	mux2_1 _RF_data_in_reg_14_U4 ( .x(n11), .d0(ALU_result[14]), .sl(mem_to_reg_EX),
		.d1(DM_read_data[14]) );
	mux2_1 _RF_data_in_reg_1_U4 ( .x(n13), .d0(ALU_result[1]), .sl(mem_to_reg_EX),
		.d1(DM_read_data[1]) );
	mux2_1 _RF_data_in_reg_9_U4 ( .x(n17), .d0(ALU_result[9]), .sl(mem_to_reg_EX),
		.d1(DM_read_data[9]) );
	smlatnr_1 mem_to_reg_MEM_reg__master ( .q(mem_to_reg_MEM_reg__m2s), .qb(),
		.d(n3), .sdi(n24), .se(test_se), .g(Ctrl__Regs_1__en1), .rb(n5), .glob_g(global_g1),
		.sync_sel(sync_sel) );
	mlatnr_2 mem_to_reg_MEM_reg__slave ( .q(mem_to_reg_MEM), .qb(), .d(mem_to_reg_MEM_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_0__master ( .q(reg_out_B_MEM_reg_0__m2s), .qb(),
		.d(reg_out_B_EX[0]), .sdi(mem_to_reg_MEM), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_0__slave ( .q(reg_out_B_MEM[0]), .qb(), .d(reg_out_B_MEM_reg_0__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_10__master ( .q(reg_out_B_MEM_reg_10__m2s),
		.qb(), .d(reg_out_B_EX[10]), .sdi(reg_out_B_MEM[9]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_10__slave ( .q(reg_out_B_MEM[10]), .qb(), .d(reg_out_B_MEM_reg_10__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_11__master ( .q(reg_out_B_MEM_reg_11__m2s),
		.qb(), .d(reg_out_B_EX[11]), .sdi(reg_out_B_MEM[10]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_11__slave ( .q(reg_out_B_MEM[11]), .qb(), .d(reg_out_B_MEM_reg_11__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_12__master ( .q(reg_out_B_MEM_reg_12__m2s),
		.qb(), .d(reg_out_B_EX[12]), .sdi(reg_out_B_MEM[11]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_12__slave ( .q(reg_out_B_MEM[12]), .qb(), .d(reg_out_B_MEM_reg_12__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_13__master ( .q(reg_out_B_MEM_reg_13__m2s),
		.qb(), .d(reg_out_B_EX[13]), .sdi(reg_out_B_MEM[12]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_13__slave ( .q(reg_out_B_MEM[13]), .qb(), .d(reg_out_B_MEM_reg_13__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_14__master ( .q(reg_out_B_MEM_reg_14__m2s),
		.qb(), .d(reg_out_B_EX[14]), .sdi(reg_out_B_MEM[13]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_14__slave ( .q(reg_out_B_MEM[14]), .qb(), .d(reg_out_B_MEM_reg_14__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_15__master ( .q(reg_out_B_MEM_reg_15__m2s),
		.qb(), .d(reg_out_B_EX[15]), .sdi(reg_out_B_MEM[14]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_15__slave ( .q(reg_out_B_MEM[15]), .qb(), .d(reg_out_B_MEM_reg_15__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_16__master ( .q(reg_out_B_MEM_reg_16__m2s),
		.qb(), .d(reg_out_B_EX[16]), .sdi(reg_out_B_MEM[15]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_16__slave ( .q(reg_out_B_MEM[16]), .qb(), .d(reg_out_B_MEM_reg_16__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_17__master ( .q(reg_out_B_MEM_reg_17__m2s),
		.qb(), .d(reg_out_B_EX[17]), .sdi(reg_out_B_MEM[16]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_17__slave ( .q(reg_out_B_MEM[17]), .qb(), .d(reg_out_B_MEM_reg_17__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_18__master ( .q(reg_out_B_MEM_reg_18__m2s),
		.qb(), .d(reg_out_B_EX[18]), .sdi(reg_out_B_MEM[17]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_18__slave ( .q(reg_out_B_MEM[18]), .qb(), .d(reg_out_B_MEM_reg_18__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_19__master ( .q(reg_out_B_MEM_reg_19__m2s),
		.qb(), .d(reg_out_B_EX[19]), .sdi(reg_out_B_MEM[18]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_19__slave ( .q(reg_out_B_MEM[19]), .qb(), .d(reg_out_B_MEM_reg_19__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_1__master ( .q(reg_out_B_MEM_reg_1__m2s), .qb(),
		.d(reg_out_B_EX[1]), .sdi(reg_out_B_MEM[0]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_1__slave ( .q(reg_out_B_MEM[1]), .qb(), .d(reg_out_B_MEM_reg_1__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_20__master ( .q(reg_out_B_MEM_reg_20__m2s),
		.qb(), .d(reg_out_B_EX[20]), .sdi(reg_out_B_MEM[19]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_20__slave ( .q(reg_out_B_MEM[20]), .qb(), .d(reg_out_B_MEM_reg_20__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_21__master ( .q(reg_out_B_MEM_reg_21__m2s),
		.qb(), .d(reg_out_B_EX[21]), .sdi(reg_out_B_MEM[20]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_21__slave ( .q(reg_out_B_MEM[21]), .qb(), .d(reg_out_B_MEM_reg_21__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_22__master ( .q(reg_out_B_MEM_reg_22__m2s),
		.qb(), .d(reg_out_B_EX[22]), .sdi(reg_out_B_MEM[21]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_22__slave ( .q(reg_out_B_MEM[22]), .qb(), .d(reg_out_B_MEM_reg_22__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_23__master ( .q(reg_out_B_MEM_reg_23__m2s),
		.qb(), .d(reg_out_B_EX[23]), .sdi(reg_out_B_MEM[22]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_23__slave ( .q(reg_out_B_MEM[23]), .qb(), .d(reg_out_B_MEM_reg_23__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_24__master ( .q(reg_out_B_MEM_reg_24__m2s),
		.qb(), .d(reg_out_B_EX[24]), .sdi(reg_out_B_MEM[23]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_24__slave ( .q(reg_out_B_MEM[24]), .qb(), .d(reg_out_B_MEM_reg_24__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_25__master ( .q(reg_out_B_MEM_reg_25__m2s),
		.qb(), .d(reg_out_B_EX[25]), .sdi(reg_out_B_MEM[24]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_25__slave ( .q(reg_out_B_MEM[25]), .qb(), .d(reg_out_B_MEM_reg_25__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_26__master ( .q(reg_out_B_MEM_reg_26__m2s),
		.qb(), .d(reg_out_B_EX[26]), .sdi(reg_out_B_MEM[25]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_26__slave ( .q(reg_out_B_MEM[26]), .qb(), .d(reg_out_B_MEM_reg_26__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_27__master ( .q(reg_out_B_MEM_reg_27__m2s),
		.qb(), .d(reg_out_B_EX[27]), .sdi(reg_out_B_MEM[26]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_27__slave ( .q(reg_out_B_MEM[27]), .qb(), .d(reg_out_B_MEM_reg_27__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_28__master ( .q(reg_out_B_MEM_reg_28__m2s),
		.qb(), .d(reg_out_B_EX[28]), .sdi(reg_out_B_MEM[27]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_28__slave ( .q(reg_out_B_MEM[28]), .qb(), .d(reg_out_B_MEM_reg_28__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_29__master ( .q(reg_out_B_MEM_reg_29__m2s),
		.qb(), .d(reg_out_B_EX[29]), .sdi(reg_out_B_MEM[28]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_29__slave ( .q(reg_out_B_MEM[29]), .qb(), .d(reg_out_B_MEM_reg_29__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_2__master ( .q(reg_out_B_MEM_reg_2__m2s), .qb(),
		.d(reg_out_B_EX[2]), .sdi(reg_out_B_MEM[1]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_2__slave ( .q(reg_out_B_MEM[2]), .qb(), .d(reg_out_B_MEM_reg_2__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_30__master ( .q(reg_out_B_MEM_reg_30__m2s),
		.qb(), .d(reg_out_B_EX[30]), .sdi(reg_out_B_MEM[29]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_30__slave ( .q(reg_out_B_MEM[30]), .qb(), .d(reg_out_B_MEM_reg_30__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_31__master ( .q(reg_out_B_MEM_reg_31__m2s),
		.qb(), .d(reg_out_B_EX[31]), .sdi(reg_out_B_MEM[30]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_31__slave ( .q(reg_out_B_MEM[31]), .qb(), .d(reg_out_B_MEM_reg_31__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_3__master ( .q(reg_out_B_MEM_reg_3__m2s), .qb(),
		.d(reg_out_B_EX[3]), .sdi(reg_out_B_MEM[2]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_3__slave ( .q(reg_out_B_MEM[3]), .qb(), .d(reg_out_B_MEM_reg_3__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_4__master ( .q(reg_out_B_MEM_reg_4__m2s), .qb(),
		.d(reg_out_B_EX[4]), .sdi(reg_out_B_MEM[3]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_4__slave ( .q(reg_out_B_MEM[4]), .qb(), .d(reg_out_B_MEM_reg_4__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_5__master ( .q(reg_out_B_MEM_reg_5__m2s), .qb(),
		.d(reg_out_B_EX[5]), .sdi(reg_out_B_MEM[4]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_5__slave ( .q(reg_out_B_MEM[5]), .qb(), .d(reg_out_B_MEM_reg_5__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_6__master ( .q(reg_out_B_MEM_reg_6__m2s), .qb(),
		.d(reg_out_B_EX[6]), .sdi(reg_out_B_MEM[5]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n5), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_6__slave ( .q(reg_out_B_MEM[6]), .qb(), .d(reg_out_B_MEM_reg_6__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n5), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_7__master ( .q(reg_out_B_MEM_reg_7__m2s), .qb(),
		.d(reg_out_B_EX[7]), .sdi(reg_out_B_MEM[6]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n4), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_7__slave ( .q(reg_out_B_MEM[7]), .qb(), .d(reg_out_B_MEM_reg_7__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n4), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_8__master ( .q(reg_out_B_MEM_reg_8__m2s), .qb(),
		.d(reg_out_B_EX[8]), .sdi(reg_out_B_MEM[7]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_8__slave ( .q(reg_out_B_MEM[8]), .qb(), .d(reg_out_B_MEM_reg_8__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_out_B_MEM_reg_9__master ( .q(reg_out_B_MEM_reg_9__m2s), .qb(),
		.d(reg_out_B_EX[9]), .sdi(reg_out_B_MEM[8]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_out_B_MEM_reg_9__slave ( .q(reg_out_B_MEM[9]), .qb(), .d(reg_out_B_MEM_reg_9__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );
	smlatnr_1 reg_write_MEM_reg__master ( .q(reg_write_MEM_reg__m2s), .qb(),
		.d(reg_write_EX), .sdi(reg_out_B_MEM[31]), .se(test_se), .g(Ctrl__Regs_1__en1),
		.rb(n6), .glob_g(global_g1), .sync_sel(sync_sel) );
	mlatnr_2 reg_write_MEM_reg__slave ( .q(reg_write_MEM), .qb(test_so), .d(reg_write_MEM_reg__m2s),
		.g(Ctrl__Regs_1__en2), .rb(n6), .glob_g(global_g2), .sync_sel(sync_sel) );

endmodule


module DLX_sync_desync (  DM_read_data, DM_write_data, DM_addr, DM_write,
	DM_read, NPC, reset, IR, byte0, word, INT, CLI, PIPEEMPTY, FREEZE, test_si,
	test_se, sync_sel, global_g1, global_g2, Ctrl__EXinst___Regs_1__en1, Ctrl__EXinst___Regs_1__en2,
	Ctrl__IDinst___Regs_1__en1, Ctrl__IDinst___Regs_1__en2, Ctrl__IFinst___Regs_1__en1,
	Ctrl__IFinst___Regs_1__en2, Ctrl__MEMinst___Regs_1__en1, Ctrl__MEMinst___Regs_1__en2 );

input  reset, INT, FREEZE, test_si, test_se, sync_sel, global_g1, global_g2,
	Ctrl__EXinst___Regs_1__en1, Ctrl__EXinst___Regs_1__en2, Ctrl__IDinst___Regs_1__en1,
	Ctrl__IDinst___Regs_1__en2, Ctrl__IFinst___Regs_1__en1, Ctrl__IFinst___Regs_1__en2,
	Ctrl__MEMinst___Regs_1__en1, Ctrl__MEMinst___Regs_1__en2;
input [31:0] DM_read_data, IR;
output  DM_write, DM_read, byte0, word, CLI, PIPEEMPTY;
output [31:0] DM_write_data, DM_addr, NPC;

wire IR_function_field_0_0, IR_function_field_1_0, IR_function_field_2_0,
	IR_function_field_3_0, IR_function_field_4_0, IR_function_field_5_0, IR_latched_0_0,
	IR_latched_10_0, IR_latched_11_0, IR_latched_12_0, IR_latched_13_0, IR_latched_14_0,
	IR_latched_15_0, IR_latched_16_0, IR_latched_17_0, IR_latched_18_0, IR_latched_19_0,
	IR_latched_1_0, IR_latched_20_0, IR_latched_21_0, IR_latched_22_0, IR_latched_23_0,
	IR_latched_24_0, IR_latched_25_0, IR_latched_26_0, IR_latched_27_0, IR_latched_28_0,
	IR_latched_29_0, IR_latched_2_0, IR_latched_30_0, IR_latched_31_0, IR_latched_3_0,
	IR_latched_4_0, IR_latched_5_0, IR_latched_6_0, IR_latched_7_0, IR_latched_8_0,
	IR_latched_9_0, IR_opcode_field_0_0, IR_opcode_field_1_0, IR_opcode_field_2_0,
	IR_opcode_field_3_0, IR_opcode_field_4_0, IR_opcode_field_5_0, Imm_0_0,
	Imm_10_0, Imm_11_0, Imm_12_0, Imm_13_0, Imm_14_0, Imm_15_0, Imm_16_0,
	Imm_17_0, Imm_18_0, Imm_19_0, Imm_1_0, Imm_20_0, Imm_21_0, Imm_22_0, Imm_23_0,
	Imm_24_0, Imm_25_0, Imm_26_0, Imm_27_0, Imm_28_0, Imm_29_0, Imm_2_0, Imm_30_0,
	Imm_31_0, Imm_3_0, Imm_4_0, Imm_5_0, Imm_6_0, Imm_7_0, Imm_8_0, Imm_9_0,
	RF_data_in_0_0, RF_data_in_10_0, RF_data_in_11_0, RF_data_in_12_0, RF_data_in_13_0,
	RF_data_in_14_0, RF_data_in_15_0, RF_data_in_16_0, RF_data_in_17_0, RF_data_in_18_0,
	RF_data_in_19_0, RF_data_in_1_0, RF_data_in_20_0, RF_data_in_21_0, RF_data_in_22_0,
	RF_data_in_23_0, RF_data_in_24_0, RF_data_in_25_0, RF_data_in_26_0, RF_data_in_27_0,
	RF_data_in_28_0, RF_data_in_29_0, RF_data_in_2_0, RF_data_in_30_0, RF_data_in_31_0,
	RF_data_in_3_0, RF_data_in_4_0, RF_data_in_5_0, RF_data_in_6_0, RF_data_in_7_0,
	RF_data_in_8_0, RF_data_in_9_0, RF_data_old_0_0, RF_data_old_10_0, RF_data_old_11_0,
	RF_data_old_12_0, RF_data_old_13_0, RF_data_old_14_0, RF_data_old_15_0,
	RF_data_old_16_0, RF_data_old_17_0, RF_data_old_18_0, RF_data_old_19_0,
	RF_data_old_1_0, RF_data_old_20_0, RF_data_old_21_0, RF_data_old_22_0,
	RF_data_old_23_0, RF_data_old_24_0, RF_data_old_25_0, RF_data_old_26_0,
	RF_data_old_27_0, RF_data_old_28_0, RF_data_old_29_0, RF_data_old_2_0,
	RF_data_old_30_0, RF_data_old_31_0, RF_data_old_3_0, RF_data_old_4_0,
	RF_data_old_5_0, RF_data_old_6_0, RF_data_old_7_0, RF_data_old_8_0, RF_data_old_9_0,
	branch_address_0_0, branch_address_10_0, branch_address_11_0, branch_address_12_0,
	branch_address_13_0, branch_address_14_0, branch_address_15_0, branch_address_16_0,
	branch_address_17_0, branch_address_18_0, branch_address_19_0, branch_address_1_0,
	branch_address_20_0, branch_address_21_0, branch_address_22_0, branch_address_23_0,
	branch_address_24_0, branch_address_25_0, branch_address_26_0, branch_address_27_0,
	branch_address_28_0, branch_address_29_0, branch_address_2_0, branch_address_30_0,
	branch_address_31_0, branch_address_3_0, branch_address_4_0, branch_address_5_0,
	branch_address_6_0, branch_address_7_0, branch_address_8_0, branch_address_9_0,
	branch_sig, counter_0_0, counter_1_0, mem_read, mem_to_reg, mem_to_reg_EX,
	mem_write, n11, n12, n13, n14, n16, n17, n2, n4, n5, n6, n8, reg_dst,
	reg_out_A_0_0, reg_out_A_10_0, reg_out_A_11_0, reg_out_A_12_0, reg_out_A_13_0,
	reg_out_A_14_0, reg_out_A_15_0, reg_out_A_16_0, reg_out_A_17_0, reg_out_A_18_0,
	reg_out_A_19_0, reg_out_A_1_0, reg_out_A_20_0, reg_out_A_21_0, reg_out_A_22_0,
	reg_out_A_23_0, reg_out_A_24_0, reg_out_A_25_0, reg_out_A_26_0, reg_out_A_27_0,
	reg_out_A_28_0, reg_out_A_29_0, reg_out_A_2_0, reg_out_A_30_0, reg_out_A_31_0,
	reg_out_A_3_0, reg_out_A_4_0, reg_out_A_5_0, reg_out_A_6_0, reg_out_A_7_0,
	reg_out_A_8_0, reg_out_A_9_0, reg_out_B_0_0, reg_out_B_10_0, reg_out_B_11_0,
	reg_out_B_12_0, reg_out_B_13_0, reg_out_B_14_0, reg_out_B_15_0, reg_out_B_16_0,
	reg_out_B_17_0, reg_out_B_18_0, reg_out_B_19_0, reg_out_B_1_0, reg_out_B_20_0,
	reg_out_B_21_0, reg_out_B_22_0, reg_out_B_23_0, reg_out_B_24_0, reg_out_B_25_0,
	reg_out_B_26_0, reg_out_B_27_0, reg_out_B_28_0, reg_out_B_29_0, reg_out_B_2_0,
	reg_out_B_30_0, reg_out_B_31_0, reg_out_B_3_0, reg_out_B_4_0, reg_out_B_5_0,
	reg_out_B_6_0, reg_out_B_7_0, reg_out_B_8_0, reg_out_B_9_0, reg_write,
	reg_write_EX, reg_write_MEM, stall;


	EX_test_1_desync EXinst ( .ALU_result(DM_addr), .reg_out_B_EX(DM_write_data),
		.mem_write_EX(DM_write), .mem_read_EX(DM_read), .mem_to_reg_EX(mem_to_reg_EX),
		.reg_write_EX(reg_write_EX), .reset(reset), .IR_opcode_field({ IR_opcode_field_5_0,
		IR_opcode_field_4_0, IR_opcode_field_3_0, IR_opcode_field_2_0, IR_opcode_field_1_0,
		IR_opcode_field_0_0}), .IR_function_field({ IR_function_field_5_0, IR_function_field_4_0,
		IR_function_field_3_0, IR_function_field_2_0, IR_function_field_1_0,
		IR_function_field_0_0}), .reg_out_A({ reg_out_A_31_0, reg_out_A_30_0,
		reg_out_A_29_0, reg_out_A_28_0, reg_out_A_27_0, reg_out_A_26_0, reg_out_A_25_0,
		reg_out_A_24_0, reg_out_A_23_0, reg_out_A_22_0, reg_out_A_21_0, reg_out_A_20_0,
		reg_out_A_19_0, reg_out_A_18_0, reg_out_A_17_0, reg_out_A_16_0, reg_out_A_15_0,
		reg_out_A_14_0, reg_out_A_13_0, reg_out_A_12_0, reg_out_A_11_0, reg_out_A_10_0,
		reg_out_A_9_0, reg_out_A_8_0, reg_out_A_7_0, reg_out_A_6_0, reg_out_A_5_0,
		reg_out_A_4_0, reg_out_A_3_0, reg_out_A_2_0, reg_out_A_1_0, reg_out_A_0_0}),
		.reg_out_B({ reg_out_B_31_0, reg_out_B_30_0, reg_out_B_29_0, reg_out_B_28_0,
		reg_out_B_27_0, reg_out_B_26_0, reg_out_B_25_0, reg_out_B_24_0, reg_out_B_23_0,
		reg_out_B_22_0, reg_out_B_21_0, reg_out_B_20_0, reg_out_B_19_0, reg_out_B_18_0,
		reg_out_B_17_0, reg_out_B_16_0, reg_out_B_15_0, reg_out_B_14_0, reg_out_B_13_0,
		reg_out_B_12_0, reg_out_B_11_0, reg_out_B_10_0, reg_out_B_9_0, reg_out_B_8_0,
		reg_out_B_7_0, reg_out_B_6_0, reg_out_B_5_0, reg_out_B_4_0, reg_out_B_3_0,
		reg_out_B_2_0, reg_out_B_1_0, reg_out_B_0_0}), .Imm({ Imm_31_0, Imm_30_0,
		Imm_29_0, Imm_28_0, Imm_27_0, Imm_26_0, Imm_25_0, Imm_24_0, Imm_23_0,
		Imm_22_0, Imm_21_0, Imm_20_0, Imm_19_0, Imm_18_0, Imm_17_0, Imm_16_0,
		Imm_15_0, Imm_14_0, Imm_13_0, Imm_12_0, Imm_11_0, Imm_10_0, Imm_9_0,
		Imm_8_0, Imm_7_0, Imm_6_0, Imm_5_0, Imm_4_0, Imm_3_0, Imm_2_0, Imm_1_0,
		Imm_0_0}), .reg_dst(reg_dst), .reg_write(reg_write), .mem_to_reg(mem_to_reg),
		.mem_read(mem_read), .mem_write(mem_write), ._byte(byte0), .word(word),
		.counter({ counter_1_0, counter_0_0}), .test_si(test_si), .test_so(n14),
		.test_se(test_se), .sync_sel(sync_sel), .global_g1(global_g1), .global_g2(global_g2),
		.Ctrl__Regs_1__en1(Ctrl__EXinst___Regs_1__en1), .Ctrl__Regs_1__en2(Ctrl__EXinst___Regs_1__en2) );
	ID_test_1_desync IDinst ( .INT(INT), .CLI(CLI), .PIPEEMPTY(PIPEEMPTY),
		.FREEZE(FREEZE), .branch_address({ branch_address_31_0, branch_address_30_0,
		branch_address_29_0, branch_address_28_0, branch_address_27_0, branch_address_26_0,
		branch_address_25_0, branch_address_24_0, branch_address_23_0, branch_address_22_0,
		branch_address_21_0, branch_address_20_0, branch_address_19_0, branch_address_18_0,
		branch_address_17_0, branch_address_16_0, branch_address_15_0, branch_address_14_0,
		branch_address_13_0, branch_address_12_0, branch_address_11_0, branch_address_10_0,
		branch_address_9_0, branch_address_8_0, branch_address_7_0, branch_address_6_0,
		branch_address_5_0, branch_address_4_0, branch_address_3_0, branch_address_2_0,
		branch_address_1_0, branch_address_0_0}), .branch_sig(branch_sig), .Imm({
		Imm_31_0, Imm_30_0, Imm_29_0, Imm_28_0, Imm_27_0, Imm_26_0, Imm_25_0,
		Imm_24_0, Imm_23_0, Imm_22_0, Imm_21_0, Imm_20_0, Imm_19_0, Imm_18_0,
		Imm_17_0, Imm_16_0, Imm_15_0, Imm_14_0, Imm_13_0, Imm_12_0, Imm_11_0,
		Imm_10_0, Imm_9_0, Imm_8_0, Imm_7_0, Imm_6_0, Imm_5_0, Imm_4_0, Imm_3_0,
		Imm_2_0, Imm_1_0, Imm_0_0}), .rt_addr(), .rd_addr(), .reg_dst(reg_dst),
		.reg_write(reg_write), .mem_to_reg(mem_to_reg), .mem_write(mem_write),
		.mem_read(mem_read), .IR_opcode_field({ IR_opcode_field_5_0, IR_opcode_field_4_0,
		IR_opcode_field_3_0, IR_opcode_field_2_0, IR_opcode_field_1_0, IR_opcode_field_0_0}),
		.IR_function_field({ IR_function_field_5_0, IR_function_field_4_0, IR_function_field_3_0,
		IR_function_field_2_0, IR_function_field_1_0, IR_function_field_0_0}),
		.stall(stall), .counter({ counter_1_0, counter_0_0}), .reset(reset),
		.NPC({ NPC[31], NPC[30], NPC[29], NPC[28], NPC[27], NPC[26], NPC[25],
		NPC[24], NPC[23], NPC[22], NPC[21], NPC[20], NPC[19], NPC[18], NPC[17],
		NPC[16], NPC[15], NPC[14], NPC[13], NPC[12], NPC[11], NPC[10], NPC[9],
		NPC[8], NPC[7], NPC[6], NPC[5], NPC[4], NPC[3], n5, NPC[1], NPC[0]}),
		.IR_latched_input({ IR_latched_31_0, IR_latched_30_0, IR_latched_29_0,
		IR_latched_28_0, IR_latched_27_0, IR_latched_26_0, IR_latched_25_0, IR_latched_24_0,
		IR_latched_23_0, IR_latched_22_0, IR_latched_21_0, IR_latched_20_0, IR_latched_19_0,
		IR_latched_18_0, IR_latched_17_0, IR_latched_16_0, IR_latched_15_0, IR_latched_14_0,
		IR_latched_13_0, IR_latched_12_0, IR_latched_11_0, IR_latched_10_0, IR_latched_9_0,
		IR_latched_8_0, IR_latched_7_0, IR_latched_6_0, IR_latched_5_0, IR_latched_4_0,
		IR_latched_3_0, IR_latched_2_0, IR_latched_1_0, IR_latched_0_0}), .reg_out_A({
		reg_out_A_31_0, reg_out_A_30_0, reg_out_A_29_0, reg_out_A_28_0, reg_out_A_27_0,
		reg_out_A_26_0, reg_out_A_25_0, reg_out_A_24_0, reg_out_A_23_0, reg_out_A_22_0,
		reg_out_A_21_0, reg_out_A_20_0, reg_out_A_19_0, reg_out_A_18_0, reg_out_A_17_0,
		reg_out_A_16_0, reg_out_A_15_0, reg_out_A_14_0, reg_out_A_13_0, reg_out_A_12_0,
		reg_out_A_11_0, reg_out_A_10_0, reg_out_A_9_0, reg_out_A_8_0, reg_out_A_7_0,
		reg_out_A_6_0, reg_out_A_5_0, reg_out_A_4_0, reg_out_A_3_0, reg_out_A_2_0,
		reg_out_A_1_0, reg_out_A_0_0}), .reg_out_B({ reg_out_B_31_0, reg_out_B_30_0,
		reg_out_B_29_0, reg_out_B_28_0, reg_out_B_27_0, reg_out_B_26_0, reg_out_B_25_0,
		reg_out_B_24_0, reg_out_B_23_0, reg_out_B_22_0, reg_out_B_21_0, reg_out_B_20_0,
		reg_out_B_19_0, reg_out_B_18_0, reg_out_B_17_0, reg_out_B_16_0, reg_out_B_15_0,
		reg_out_B_14_0, reg_out_B_13_0, reg_out_B_12_0, reg_out_B_11_0, reg_out_B_10_0,
		reg_out_B_9_0, reg_out_B_8_0, reg_out_B_7_0, reg_out_B_6_0, reg_out_B_5_0,
		reg_out_B_4_0, reg_out_B_3_0, reg_out_B_2_0, reg_out_B_1_0, reg_out_B_0_0}),
		.reg_write_WB(reg_write_MEM), .WB_data({ RF_data_in_31_0, RF_data_in_30_0,
		RF_data_in_29_0, RF_data_in_28_0, RF_data_in_27_0, RF_data_in_26_0, RF_data_in_25_0,
		RF_data_in_24_0, RF_data_in_23_0, RF_data_in_22_0, RF_data_in_21_0, RF_data_in_20_0,
		RF_data_in_19_0, RF_data_in_18_0, RF_data_in_17_0, RF_data_in_16_0, RF_data_in_15_0,
		RF_data_in_14_0, RF_data_in_13_0, RF_data_in_12_0, RF_data_in_11_0, RF_data_in_10_0,
		RF_data_in_9_0, RF_data_in_8_0, RF_data_in_7_0, RF_data_in_6_0, RF_data_in_5_0,
		RF_data_in_4_0, RF_data_in_3_0, RF_data_in_2_0, RF_data_in_1_0, RF_data_in_0_0}),
		.WB_data_old({ RF_data_old_31_0, RF_data_old_30_0, RF_data_old_29_0,
		RF_data_old_28_0, RF_data_old_27_0, RF_data_old_26_0, RF_data_old_25_0,
		RF_data_old_24_0, RF_data_old_23_0, RF_data_old_22_0, RF_data_old_21_0,
		RF_data_old_20_0, RF_data_old_19_0, RF_data_old_18_0, RF_data_old_17_0,
		RF_data_old_16_0, RF_data_old_15_0, RF_data_old_14_0, RF_data_old_13_0,
		RF_data_old_12_0, RF_data_old_11_0, RF_data_old_10_0, RF_data_old_9_0,
		RF_data_old_8_0, RF_data_old_7_0, RF_data_old_6_0, RF_data_old_5_0, RF_data_old_4_0,
		RF_data_old_3_0, RF_data_old_2_0, RF_data_old_1_0, RF_data_old_0_0}),
		.test_si(n14), .test_so(n13), .test_se(test_se), .sync_sel(sync_sel),
		.global_g1(global_g1), .global_g2(global_g2), .Ctrl__Regs_1__en1(Ctrl__IDinst___Regs_1__en1),
		.Ctrl__Regs_1__en2(Ctrl__IDinst___Regs_1__en2) );
	IF_test_1_desync IFinst ( .NPC({ NPC[31], NPC[30], NPC[29], NPC[28], NPC[27],
		NPC[26], NPC[25], NPC[24], NPC[23], NPC[22], NPC[21], NPC[20], NPC[19],
		NPC[18], NPC[17], NPC[16], NPC[15], NPC[14], NPC[13], n4, NPC[11], n16,
		NPC[9], NPC[8], n17, NPC[6], NPC[5], NPC[4], NPC[3], n5, NPC[1], NPC[0]}),
		.PC(), .IR_latched({ IR_latched_31_0, IR_latched_30_0, IR_latched_29_0,
		IR_latched_28_0, IR_latched_27_0, IR_latched_26_0, IR_latched_25_0, IR_latched_24_0,
		IR_latched_23_0, IR_latched_22_0, IR_latched_21_0, IR_latched_20_0, IR_latched_19_0,
		IR_latched_18_0, IR_latched_17_0, IR_latched_16_0, IR_latched_15_0, IR_latched_14_0,
		IR_latched_13_0, IR_latched_12_0, IR_latched_11_0, IR_latched_10_0, IR_latched_9_0,
		IR_latched_8_0, IR_latched_7_0, IR_latched_6_0, IR_latched_5_0, IR_latched_4_0,
		IR_latched_3_0, IR_latched_2_0, IR_latched_1_0, IR_latched_0_0}), .reset(reset),
		.branch_sig(branch_sig), .branch_address({ branch_address_31_0, branch_address_30_0,
		branch_address_29_0, branch_address_28_0, branch_address_27_0, branch_address_26_0,
		branch_address_25_0, branch_address_24_0, branch_address_23_0, branch_address_22_0,
		branch_address_21_0, branch_address_20_0, branch_address_19_0, branch_address_18_0,
		branch_address_17_0, branch_address_16_0, branch_address_15_0, branch_address_14_0,
		branch_address_13_0, branch_address_12_0, branch_address_11_0, branch_address_10_0,
		branch_address_9_0, branch_address_8_0, branch_address_7_0, branch_address_6_0,
		branch_address_5_0, branch_address_4_0, branch_address_3_0, branch_address_2_0,
		branch_address_1_0, branch_address_0_0}), .IR(IR), .stall(stall), .counter({
		counter_1_0, counter_0_0}), .test_si1(n13), .test_so1(n12), .test_si2(n11),
		.test_se(test_se), .sync_sel(sync_sel), .global_g1(global_g1), .global_g2(global_g2),
		.Ctrl__Regs_1__en1(Ctrl__IFinst___Regs_1__en1), .Ctrl__Regs_1__en2(Ctrl__IFinst___Regs_1__en2) );
	MEM_test_1_desync MEMinst ( .reg_write_MEM(reg_write_MEM), .mem_to_reg_EX(mem_to_reg_EX),
		.reset(reset), .ALU_result(DM_addr), .reg_write_EX(reg_write_EX), .mem_to_reg_MEM(),
		.reg_out_B_EX(DM_write_data), .reg_out_B_MEM({ RF_data_old_31_0, RF_data_old_30_0,
		RF_data_old_29_0, RF_data_old_28_0, RF_data_old_27_0, RF_data_old_26_0,
		RF_data_old_25_0, RF_data_old_24_0, RF_data_old_23_0, RF_data_old_22_0,
		RF_data_old_21_0, RF_data_old_20_0, RF_data_old_19_0, RF_data_old_18_0,
		RF_data_old_17_0, RF_data_old_16_0, RF_data_old_15_0, RF_data_old_14_0,
		RF_data_old_13_0, RF_data_old_12_0, RF_data_old_11_0, RF_data_old_10_0,
		RF_data_old_9_0, RF_data_old_8_0, RF_data_old_7_0, RF_data_old_6_0, RF_data_old_5_0,
		RF_data_old_4_0, RF_data_old_3_0, RF_data_old_2_0, RF_data_old_1_0, RF_data_old_0_0}),
		.DM_read_data(DM_read_data), .RF_data_in({ RF_data_in_31_0, RF_data_in_30_0,
		RF_data_in_29_0, RF_data_in_28_0, RF_data_in_27_0, RF_data_in_26_0, RF_data_in_25_0,
		RF_data_in_24_0, RF_data_in_23_0, RF_data_in_22_0, RF_data_in_21_0, RF_data_in_20_0,
		RF_data_in_19_0, RF_data_in_18_0, RF_data_in_17_0, RF_data_in_16_0, RF_data_in_15_0,
		RF_data_in_14_0, RF_data_in_13_0, RF_data_in_12_0, RF_data_in_11_0, RF_data_in_10_0,
		RF_data_in_9_0, RF_data_in_8_0, RF_data_in_7_0, RF_data_in_6_0, RF_data_in_5_0,
		RF_data_in_4_0, RF_data_in_3_0, RF_data_in_2_0, RF_data_in_1_0, RF_data_in_0_0}),
		.test_si(n12), .test_so(n11), .test_se(test_se), .sync_sel(sync_sel),
		.global_g1(global_g1), .global_g2(global_g2), .Ctrl__Regs_1__en1(Ctrl__MEMinst___Regs_1__en1),
		.Ctrl__Regs_1__en2(Ctrl__MEMinst___Regs_1__en2) );
	buf_10 U1 ( .x(NPC[12]), .a(n4) );
	inv_0 U2 ( .x(n2), .a(n5) );
	inv_2 U3 ( .x(NPC[2]), .a(n2) );
	inv_6 U4 ( .x(n6), .a(n16) );
	inv_10 U5 ( .x(NPC[10]), .a(n6) );
	inv_6 U6 ( .x(n8), .a(n17) );
	inv_10 U7 ( .x(NPC[7]), .a(n8) );

endmodule


module DLX_sync_desync_with_ctrls (  DM_read_data, DM_write_data, DM_addr,
	DM_write, DM_read, NPC, reset, IR, byte0, word, INT, CLI, PIPEEMPTY, FREEZE,
	test_si, test_se, sync_sel, global_g1, global_g2, Ctrl__reset, Ctrl__EXinst___Regs_1__ai,
	Ctrl__IDinst___Regs_1__ai, Ctrl__IDinst___Regs_1__ro, Ctrl__MEMinst___Regs_1__ro,
	Ctrl__IFinst___Regs_1__ri, Ctrl__IFinst___Regs_1__ai, Ctrl__MEMinst___Regs_1__ri,
	Ctrl__MEMinst___Regs_1__ai, Ctrl__EXinst___Regs_1__ro, Ctrl__EXinst___Regs_1__ao,
	Ctrl__IFinst___Regs_1__ro, Ctrl__IFinst___Regs_1__ao, Ctrl__EXinst___Regs_1__delay_mux_sel,
	Ctrl__IDinst___Regs_1__delay_mux_sel, Ctrl__IFinst___Regs_1__delay_mux_sel,
	Ctrl__MEMinst___Regs_1__delay_mux_sel, Ctrl__EXinst___Regs_1__en1, Ctrl__EXinst___Regs_1__en2,
	Ctrl__IDinst___Regs_1__en1, Ctrl__IDinst___Regs_1__en2, Ctrl__IFinst___Regs_1__en1,
	Ctrl__IFinst___Regs_1__en2, Ctrl__MEMinst___Regs_1__en1, Ctrl__MEMinst___Regs_1__en2/*,
	Ctrl__EXinst___Regs_1__en1_new, Ctrl__EXinst___Regs_1__en2_new, Ctrl__IFinst___Regs_1__en1_new,
	Ctrl__IFinst___Regs_1__en2_new, Ctrl__IDinst___Regs_1__en1_new, Ctrl__IDinst___Regs_1__en2_new,
	Ctrl__MEMinst___Regs_1__en1_new, Ctrl__MEMinst___Regs_1__en2_new*/ );

input  reset, INT, FREEZE, test_si, test_se, sync_sel, global_g1, global_g2,
	Ctrl__reset, Ctrl__IFinst___Regs_1__ri, Ctrl__MEMinst___Regs_1__ri,
	Ctrl__EXinst___Regs_1__ao, Ctrl__IFinst___Regs_1__ao/*, Ctrl__EXinst___Regs_1__en1_new,
	Ctrl__EXinst___Regs_1__en2_new, Ctrl__IFinst___Regs_1__en1_new, Ctrl__IFinst___Regs_1__en2_new,
	Ctrl__IDinst___Regs_1__en1_new, Ctrl__IDinst___Regs_1__en2_new, Ctrl__MEMinst___Regs_1__en1_new,
	Ctrl__MEMinst___Regs_1__en2_new*/;
input [1:0] Ctrl__EXinst___Regs_1__delay_mux_sel, Ctrl__IDinst___Regs_1__delay_mux_sel,
	Ctrl__IFinst___Regs_1__delay_mux_sel, Ctrl__MEMinst___Regs_1__delay_mux_sel;
input [31:0] DM_read_data, IR;
output  DM_write, DM_read, byte0, word, CLI, PIPEEMPTY, Ctrl__IDinst___Regs_1__ai,
	Ctrl__EXinst___Regs_1__ai, Ctrl__IDinst___Regs_1__ro, Ctrl__MEMinst___Regs_1__ro,
        Ctrl__IFinst___Regs_1__ai, Ctrl__MEMinst___Regs_1__ai, Ctrl__EXinst___Regs_1__ro,
        Ctrl__IFinst___Regs_1__ro, Ctrl__EXinst___Regs_1__en1, Ctrl__EXinst___Regs_1__en2,
	Ctrl__IDinst___Regs_1__en1, Ctrl__IDinst___Regs_1__en2, Ctrl__IFinst___Regs_1__en1,
	Ctrl__IFinst___Regs_1__en2, Ctrl__MEMinst___Regs_1__en1, Ctrl__MEMinst___Regs_1__en2;
output [31:0] DM_write_data, DM_addr, NPC;


	controller_d32__0_85__1__1_38__1_77_r1_a2 Ctrl__EXinst___Regs_1 ( .reset(Ctrl__reset),
		.en1(Ctrl__EXinst___Regs_1__en1), .en2(Ctrl__EXinst___Regs_1__en2), .ri1(Ctrl__IDinst___Regs_1__ro),
		.ai(Ctrl__EXinst___Regs_1__ai), .ro(Ctrl__EXinst___Regs_1__ro), .ao1(Ctrl__EXinst___Regs_1__ao),
		.ao2(Ctrl__MEMinst___Regs_1__ai), .delay_mux_sel(Ctrl__EXinst___Regs_1__delay_mux_sel) );
	controller_d31__0_85__1__1_47__1_93_r2_a2 Ctrl__IDinst___Regs_1 ( .reset(Ctrl__reset),
		.en1(Ctrl__IDinst___Regs_1__en1), .en2(Ctrl__IDinst___Regs_1__en2), .ri1(Ctrl__IFinst___Regs_1__ro),
		.ri2(Ctrl__MEMinst___Regs_1__ro), .ai(Ctrl__IDinst___Regs_1__ai), .ro(Ctrl__IDinst___Regs_1__ro),
		.ao1(Ctrl__EXinst___Regs_1__ai), .ao2(Ctrl__IFinst___Regs_1__ai), .delay_mux_sel(Ctrl__IDinst___Regs_1__delay_mux_sel) );
	controller_d28__0_85__1__1_48__1_95_r2_a2 Ctrl__IFinst___Regs_1 ( .reset(Ctrl__reset),
		.en1(Ctrl__IFinst___Regs_1__en1), .en2(Ctrl__IFinst___Regs_1__en2), .ri1(Ctrl__IFinst___Regs_1__ri),
		.ri2(Ctrl__IDinst___Regs_1__ro), .ai(Ctrl__IFinst___Regs_1__ai), .ro(Ctrl__IFinst___Regs_1__ro),
		.ao1(Ctrl__IFinst___Regs_1__ao), .ao2(Ctrl__IDinst___Regs_1__ai), .delay_mux_sel(Ctrl__IFinst___Regs_1__delay_mux_sel) );
	controller_d6__0_85__1__1_18__1_36_r2_a1 Ctrl__MEMinst___Regs_1 ( .reset(Ctrl__reset),
		.en1(Ctrl__MEMinst___Regs_1__en1), .en2(Ctrl__MEMinst___Regs_1__en2),
		.ri1(Ctrl__MEMinst___Regs_1__ri), .ri2(Ctrl__EXinst___Regs_1__ro), .ai(Ctrl__MEMinst___Regs_1__ai),
		.ro(Ctrl__MEMinst___Regs_1__ro), .ao1(Ctrl__IDinst___Regs_1__ai), .delay_mux_sel(Ctrl__MEMinst___Regs_1__delay_mux_sel) );
	DLX_sync_desync DLX_sync ( .DM_read_data(DM_read_data), .DM_write_data(DM_write_data),
		.DM_addr(DM_addr), .DM_write(DM_write), .DM_read(DM_read), .NPC(NPC),
		.reset(reset), .IR(IR), .byte0(byte0), .word(word), .INT(INT), .CLI(CLI),
		.PIPEEMPTY(PIPEEMPTY), .FREEZE(FREEZE), .test_si(test_si), .test_se(test_se),
		.sync_sel(sync_sel), .global_g1(global_g1), .global_g2(global_g2), .Ctrl__EXinst___Regs_1__en1(Ctrl__EXinst___Regs_1__en1/*new*/),
		.Ctrl__EXinst___Regs_1__en2(Ctrl__EXinst___Regs_1__en2/*new*/), .Ctrl__IDinst___Regs_1__en1(Ctrl__IDinst___Regs_1__en1/*new*/),
		.Ctrl__IDinst___Regs_1__en2(Ctrl__IDinst___Regs_1__en2/*new*/), .Ctrl__IFinst___Regs_1__en1(Ctrl__IFinst___Regs_1__en1/*new*/),
		.Ctrl__IFinst___Regs_1__en2(Ctrl__IFinst___Regs_1__en2/*new*/), .Ctrl__MEMinst___Regs_1__en1(Ctrl__MEMinst___Regs_1__en1/*new*/),
		.Ctrl__MEMinst___Regs_1__en2(Ctrl__MEMinst___Regs_1__en2/*new*/) );

endmodule


