module abc (id3, id4);
    input id3;
    output id4;

    a = vector1[5] + vector[6];
    b = vector2[WIDTH] + vector3[6];
    c = vector3[4:6] + vectro4[5] + vector[WIDTH];
    d = vector5[6 +: WIDTH];
    f = vector5[WIDTH -: 5];
    g = vector6[4 +: functionr(2134)];
    h = vector6[4 -: functionr(2134)];

    $write("a = %b, %b",id3,id4);

endmodule
