module abc (id3, id4);
    input id3;
    output id4;
    function automatic [63:0] factorial (input reg [31:0] n,t,r,input [31:0] w,c);
        a = 2;
    endfunction

    function real multiply;
        input a, b;
        real v,c;
        real a;
        a = 2;
    endfunction

    function real multiply;
        input a, b;
        a = 2;
    endfunction

    function Parity_Calc_Func;
         input [31:0] addr;
         input [31:0] addr2;
         real v,c;
         a = 2;
    endfunction

    function automatic Parity_Calc_Func;
         input [31:0] addr;
         real v,c;
         a = 2;
    endfunction

endmodule
